module top (
    input wire clk,
    input wire [30:0] io_in,
    output wire [30:0] io_out,
    io_oeb,
    output wire [7:0] bram0_rd_addr,
    bram0_wr_addr,
    output wire [31:0] bram0_wr_data,
    input wire [31:0] bram0_rd_data,
    output wire [7:0] bram0_config,
    output wire [7:0] bram1_rd_addr,
    bram1_wr_addr,
    output wire [31:0] bram1_wr_data,
    input wire [31:0] bram1_rd_data,
    output wire [7:0] bram1_config,
    output wire [7:0] bram2_rd_addr,
    bram2_wr_addr,
    output wire [31:0] bram2_wr_data,
    input wire [31:0] bram2_rd_data,
    output wire [7:0] bram2_config,
    output wire [7:0] bram3_rd_addr,
    bram3_wr_addr,
    output wire [31:0] bram3_wr_data,
    input wire [31:0] bram3_rd_data,
    output wire [7:0] bram3_config,
    output wire [7:0] bram4_rd_addr,
    bram4_wr_addr,
    output wire [31:0] bram4_wr_data,
    input wire [31:0] bram4_rd_data,
    output wire [7:0] bram4_config,
    output wire [7:0] bram5_rd_addr,
    bram5_wr_addr,
    output wire [31:0] bram5_wr_data,
    input wire [31:0] bram5_rd_data,
    output wire [7:0] bram5_config,
    output wire [7:0] bram6_rd_addr,
    bram6_wr_addr,
    output wire [31:0] bram6_wr_data,
    input wire [31:0] bram6_rd_data,
    output wire [7:0] bram6_config,
    output wire [7:0] bram7_rd_addr,
    bram7_wr_addr,
    output wire [31:0] bram7_wr_data,
    input wire [31:0] bram7_rd_data,
    output wire [7:0] bram7_config
);
    localparam N = 893;
    wire [N:0] osc;
    genvar ii;
    generate
        for (ii = 0; ii < N; ii = ii + 1'b1) begin
            LUT4 #(
                .INIT(16'h00FF)
            ) l0 (
                .I3(osc[ii]),
                .O (osc[ii+1'b1])
            );
        end
    endgenerate

    assign osc[0] = osc[N];

    wire osco;
    LUT1 #(
        .INIT(2'b1)
    ) lo (
        .I0(osc[0]),
        .O (osco)
    );

    assign io_out[23] = osco;
    assign io_oeb = ~(28'b1);
endmodule
