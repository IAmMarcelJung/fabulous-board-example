//NumberOfConfigBits:412
module RegFile_switch_matrix (
    N1END0,
    N1END1,
    N1END2,
    N1END3,
    N2MID0,
    N2MID1,
    N2MID2,
    N2MID3,
    N2MID4,
    N2MID5,
    N2MID6,
    N2MID7,
    N2END0,
    N2END1,
    N2END2,
    N2END3,
    N2END4,
    N2END5,
    N2END6,
    N2END7,
    N4END0,
    N4END1,
    N4END2,
    N4END3,
    NN4END0,
    NN4END1,
    NN4END2,
    NN4END3,
    E1END0,
    E1END1,
    E1END2,
    E1END3,
    E2MID0,
    E2MID1,
    E2MID2,
    E2MID3,
    E2MID4,
    E2MID5,
    E2MID6,
    E2MID7,
    E2END0,
    E2END1,
    E2END2,
    E2END3,
    E2END4,
    E2END5,
    E2END6,
    E2END7,
    EE4END0,
    EE4END1,
    EE4END2,
    EE4END3,
    E6END0,
    E6END1,
    S1END0,
    S1END1,
    S1END2,
    S1END3,
    S2MID0,
    S2MID1,
    S2MID2,
    S2MID3,
    S2MID4,
    S2MID5,
    S2MID6,
    S2MID7,
    S2END0,
    S2END1,
    S2END2,
    S2END3,
    S2END4,
    S2END5,
    S2END6,
    S2END7,
    S4END0,
    S4END1,
    S4END2,
    S4END3,
    SS4END0,
    SS4END1,
    SS4END2,
    SS4END3,
    W1END0,
    W1END1,
    W1END2,
    W1END3,
    W2MID0,
    W2MID1,
    W2MID2,
    W2MID3,
    W2MID4,
    W2MID5,
    W2MID6,
    W2MID7,
    W2END0,
    W2END1,
    W2END2,
    W2END3,
    W2END4,
    W2END5,
    W2END6,
    W2END7,
    WW4END0,
    WW4END1,
    WW4END2,
    WW4END3,
    W6END0,
    W6END1,
    AD0,
    AD1,
    AD2,
    AD3,
    BD0,
    BD1,
    BD2,
    BD3,
    J2MID_ABa_END0,
    J2MID_ABa_END1,
    J2MID_ABa_END2,
    J2MID_ABa_END3,
    J2MID_CDa_END0,
    J2MID_CDa_END1,
    J2MID_CDa_END2,
    J2MID_CDa_END3,
    J2MID_EFa_END0,
    J2MID_EFa_END1,
    J2MID_EFa_END2,
    J2MID_EFa_END3,
    J2MID_GHa_END0,
    J2MID_GHa_END1,
    J2MID_GHa_END2,
    J2MID_GHa_END3,
    J2MID_ABb_END0,
    J2MID_ABb_END1,
    J2MID_ABb_END2,
    J2MID_ABb_END3,
    J2MID_CDb_END0,
    J2MID_CDb_END1,
    J2MID_CDb_END2,
    J2MID_CDb_END3,
    J2MID_EFb_END0,
    J2MID_EFb_END1,
    J2MID_EFb_END2,
    J2MID_EFb_END3,
    J2MID_GHb_END0,
    J2MID_GHb_END1,
    J2MID_GHb_END2,
    J2MID_GHb_END3,
    J2END_AB_END0,
    J2END_AB_END1,
    J2END_AB_END2,
    J2END_AB_END3,
    J2END_CD_END0,
    J2END_CD_END1,
    J2END_CD_END2,
    J2END_CD_END3,
    J2END_EF_END0,
    J2END_EF_END1,
    J2END_EF_END2,
    J2END_EF_END3,
    J2END_GH_END0,
    J2END_GH_END1,
    J2END_GH_END2,
    J2END_GH_END3,
    JN2END0,
    JN2END1,
    JN2END2,
    JN2END3,
    JN2END4,
    JN2END5,
    JN2END6,
    JN2END7,
    JE2END0,
    JE2END1,
    JE2END2,
    JE2END3,
    JE2END4,
    JE2END5,
    JE2END6,
    JE2END7,
    JS2END0,
    JS2END1,
    JS2END2,
    JS2END3,
    JS2END4,
    JS2END5,
    JS2END6,
    JS2END7,
    JW2END0,
    JW2END1,
    JW2END2,
    JW2END3,
    JW2END4,
    JW2END5,
    JW2END6,
    JW2END7,
    J_l_AB_END0,
    J_l_AB_END1,
    J_l_AB_END2,
    J_l_AB_END3,
    J_l_CD_END0,
    J_l_CD_END1,
    J_l_CD_END2,
    J_l_CD_END3,
    J_l_EF_END0,
    J_l_EF_END1,
    J_l_EF_END2,
    J_l_EF_END3,
    J_l_GH_END0,
    J_l_GH_END1,
    J_l_GH_END2,
    J_l_GH_END3,
    N1BEG0,
    N1BEG1,
    N1BEG2,
    N1BEG3,
    N2BEG0,
    N2BEG1,
    N2BEG2,
    N2BEG3,
    N2BEG4,
    N2BEG5,
    N2BEG6,
    N2BEG7,
    N2BEGb0,
    N2BEGb1,
    N2BEGb2,
    N2BEGb3,
    N2BEGb4,
    N2BEGb5,
    N2BEGb6,
    N2BEGb7,
    N4BEG0,
    N4BEG1,
    N4BEG2,
    N4BEG3,
    NN4BEG0,
    NN4BEG1,
    NN4BEG2,
    NN4BEG3,
    E1BEG0,
    E1BEG1,
    E1BEG2,
    E1BEG3,
    E2BEG0,
    E2BEG1,
    E2BEG2,
    E2BEG3,
    E2BEG4,
    E2BEG5,
    E2BEG6,
    E2BEG7,
    E2BEGb0,
    E2BEGb1,
    E2BEGb2,
    E2BEGb3,
    E2BEGb4,
    E2BEGb5,
    E2BEGb6,
    E2BEGb7,
    EE4BEG0,
    EE4BEG1,
    EE4BEG2,
    EE4BEG3,
    E6BEG0,
    E6BEG1,
    S1BEG0,
    S1BEG1,
    S1BEG2,
    S1BEG3,
    S2BEG0,
    S2BEG1,
    S2BEG2,
    S2BEG3,
    S2BEG4,
    S2BEG5,
    S2BEG6,
    S2BEG7,
    S2BEGb0,
    S2BEGb1,
    S2BEGb2,
    S2BEGb3,
    S2BEGb4,
    S2BEGb5,
    S2BEGb6,
    S2BEGb7,
    S4BEG0,
    S4BEG1,
    S4BEG2,
    S4BEG3,
    SS4BEG0,
    SS4BEG1,
    SS4BEG2,
    SS4BEG3,
    W1BEG0,
    W1BEG1,
    W1BEG2,
    W1BEG3,
    W2BEG0,
    W2BEG1,
    W2BEG2,
    W2BEG3,
    W2BEG4,
    W2BEG5,
    W2BEG6,
    W2BEG7,
    W2BEGb0,
    W2BEGb1,
    W2BEGb2,
    W2BEGb3,
    W2BEGb4,
    W2BEGb5,
    W2BEGb6,
    W2BEGb7,
    WW4BEG0,
    WW4BEG1,
    WW4BEG2,
    WW4BEG3,
    W6BEG0,
    W6BEG1,
    D0,
    D1,
    D2,
    D3,
    W_ADR0,
    W_ADR1,
    W_ADR2,
    W_ADR3,
    W_ADR4,
    W_en,
    A_ADR0,
    A_ADR1,
    A_ADR2,
    A_ADR3,
    A_ADR4,
    B_ADR0,
    B_ADR1,
    B_ADR2,
    B_ADR3,
    B_ADR4,
    J2MID_ABa_BEG0,
    J2MID_ABa_BEG1,
    J2MID_ABa_BEG2,
    J2MID_ABa_BEG3,
    J2MID_CDa_BEG0,
    J2MID_CDa_BEG1,
    J2MID_CDa_BEG2,
    J2MID_CDa_BEG3,
    J2MID_EFa_BEG0,
    J2MID_EFa_BEG1,
    J2MID_EFa_BEG2,
    J2MID_EFa_BEG3,
    J2MID_GHa_BEG0,
    J2MID_GHa_BEG1,
    J2MID_GHa_BEG2,
    J2MID_GHa_BEG3,
    J2MID_ABb_BEG0,
    J2MID_ABb_BEG1,
    J2MID_ABb_BEG2,
    J2MID_ABb_BEG3,
    J2MID_CDb_BEG0,
    J2MID_CDb_BEG1,
    J2MID_CDb_BEG2,
    J2MID_CDb_BEG3,
    J2MID_EFb_BEG0,
    J2MID_EFb_BEG1,
    J2MID_EFb_BEG2,
    J2MID_EFb_BEG3,
    J2MID_GHb_BEG0,
    J2MID_GHb_BEG1,
    J2MID_GHb_BEG2,
    J2MID_GHb_BEG3,
    J2END_AB_BEG0,
    J2END_AB_BEG1,
    J2END_AB_BEG2,
    J2END_AB_BEG3,
    J2END_CD_BEG0,
    J2END_CD_BEG1,
    J2END_CD_BEG2,
    J2END_CD_BEG3,
    J2END_EF_BEG0,
    J2END_EF_BEG1,
    J2END_EF_BEG2,
    J2END_EF_BEG3,
    J2END_GH_BEG0,
    J2END_GH_BEG1,
    J2END_GH_BEG2,
    J2END_GH_BEG3,
    JN2BEG0,
    JN2BEG1,
    JN2BEG2,
    JN2BEG3,
    JN2BEG4,
    JN2BEG5,
    JN2BEG6,
    JN2BEG7,
    JE2BEG0,
    JE2BEG1,
    JE2BEG2,
    JE2BEG3,
    JE2BEG4,
    JE2BEG5,
    JE2BEG6,
    JE2BEG7,
    JS2BEG0,
    JS2BEG1,
    JS2BEG2,
    JS2BEG3,
    JS2BEG4,
    JS2BEG5,
    JS2BEG6,
    JS2BEG7,
    JW2BEG0,
    JW2BEG1,
    JW2BEG2,
    JW2BEG3,
    JW2BEG4,
    JW2BEG5,
    JW2BEG6,
    JW2BEG7,
    J_l_AB_BEG0,
    J_l_AB_BEG1,
    J_l_AB_BEG2,
    J_l_AB_BEG3,
    J_l_CD_BEG0,
    J_l_CD_BEG1,
    J_l_CD_BEG2,
    J_l_CD_BEG3,
    J_l_EF_BEG0,
    J_l_EF_BEG1,
    J_l_EF_BEG2,
    J_l_EF_BEG3,
    J_l_GH_BEG0,
    J_l_GH_BEG1,
    J_l_GH_BEG2,
    J_l_GH_BEG3,
    ConfigBits,
    ConfigBits_N
);
  parameter NoConfigBits = 412;
  // switch matrix inputs
  input N1END0;
  input N1END1;
  input N1END2;
  input N1END3;
  input N2MID0;
  input N2MID1;
  input N2MID2;
  input N2MID3;
  input N2MID4;
  input N2MID5;
  input N2MID6;
  input N2MID7;
  input N2END0;
  input N2END1;
  input N2END2;
  input N2END3;
  input N2END4;
  input N2END5;
  input N2END6;
  input N2END7;
  input N4END0;
  input N4END1;
  input N4END2;
  input N4END3;
  input NN4END0;
  input NN4END1;
  input NN4END2;
  input NN4END3;
  input E1END0;
  input E1END1;
  input E1END2;
  input E1END3;
  input E2MID0;
  input E2MID1;
  input E2MID2;
  input E2MID3;
  input E2MID4;
  input E2MID5;
  input E2MID6;
  input E2MID7;
  input E2END0;
  input E2END1;
  input E2END2;
  input E2END3;
  input E2END4;
  input E2END5;
  input E2END6;
  input E2END7;
  input EE4END0;
  input EE4END1;
  input EE4END2;
  input EE4END3;
  input E6END0;
  input E6END1;
  input S1END0;
  input S1END1;
  input S1END2;
  input S1END3;
  input S2MID0;
  input S2MID1;
  input S2MID2;
  input S2MID3;
  input S2MID4;
  input S2MID5;
  input S2MID6;
  input S2MID7;
  input S2END0;
  input S2END1;
  input S2END2;
  input S2END3;
  input S2END4;
  input S2END5;
  input S2END6;
  input S2END7;
  input S4END0;
  input S4END1;
  input S4END2;
  input S4END3;
  input SS4END0;
  input SS4END1;
  input SS4END2;
  input SS4END3;
  input W1END0;
  input W1END1;
  input W1END2;
  input W1END3;
  input W2MID0;
  input W2MID1;
  input W2MID2;
  input W2MID3;
  input W2MID4;
  input W2MID5;
  input W2MID6;
  input W2MID7;
  input W2END0;
  input W2END1;
  input W2END2;
  input W2END3;
  input W2END4;
  input W2END5;
  input W2END6;
  input W2END7;
  input WW4END0;
  input WW4END1;
  input WW4END2;
  input WW4END3;
  input W6END0;
  input W6END1;
  input AD0;
  input AD1;
  input AD2;
  input AD3;
  input BD0;
  input BD1;
  input BD2;
  input BD3;
  input J2MID_ABa_END0;
  input J2MID_ABa_END1;
  input J2MID_ABa_END2;
  input J2MID_ABa_END3;
  input J2MID_CDa_END0;
  input J2MID_CDa_END1;
  input J2MID_CDa_END2;
  input J2MID_CDa_END3;
  input J2MID_EFa_END0;
  input J2MID_EFa_END1;
  input J2MID_EFa_END2;
  input J2MID_EFa_END3;
  input J2MID_GHa_END0;
  input J2MID_GHa_END1;
  input J2MID_GHa_END2;
  input J2MID_GHa_END3;
  input J2MID_ABb_END0;
  input J2MID_ABb_END1;
  input J2MID_ABb_END2;
  input J2MID_ABb_END3;
  input J2MID_CDb_END0;
  input J2MID_CDb_END1;
  input J2MID_CDb_END2;
  input J2MID_CDb_END3;
  input J2MID_EFb_END0;
  input J2MID_EFb_END1;
  input J2MID_EFb_END2;
  input J2MID_EFb_END3;
  input J2MID_GHb_END0;
  input J2MID_GHb_END1;
  input J2MID_GHb_END2;
  input J2MID_GHb_END3;
  input J2END_AB_END0;
  input J2END_AB_END1;
  input J2END_AB_END2;
  input J2END_AB_END3;
  input J2END_CD_END0;
  input J2END_CD_END1;
  input J2END_CD_END2;
  input J2END_CD_END3;
  input J2END_EF_END0;
  input J2END_EF_END1;
  input J2END_EF_END2;
  input J2END_EF_END3;
  input J2END_GH_END0;
  input J2END_GH_END1;
  input J2END_GH_END2;
  input J2END_GH_END3;
  input JN2END0;
  input JN2END1;
  input JN2END2;
  input JN2END3;
  input JN2END4;
  input JN2END5;
  input JN2END6;
  input JN2END7;
  input JE2END0;
  input JE2END1;
  input JE2END2;
  input JE2END3;
  input JE2END4;
  input JE2END5;
  input JE2END6;
  input JE2END7;
  input JS2END0;
  input JS2END1;
  input JS2END2;
  input JS2END3;
  input JS2END4;
  input JS2END5;
  input JS2END6;
  input JS2END7;
  input JW2END0;
  input JW2END1;
  input JW2END2;
  input JW2END3;
  input JW2END4;
  input JW2END5;
  input JW2END6;
  input JW2END7;
  input J_l_AB_END0;
  input J_l_AB_END1;
  input J_l_AB_END2;
  input J_l_AB_END3;
  input J_l_CD_END0;
  input J_l_CD_END1;
  input J_l_CD_END2;
  input J_l_CD_END3;
  input J_l_EF_END0;
  input J_l_EF_END1;
  input J_l_EF_END2;
  input J_l_EF_END3;
  input J_l_GH_END0;
  input J_l_GH_END1;
  input J_l_GH_END2;
  input J_l_GH_END3;
  output N1BEG0;
  output N1BEG1;
  output N1BEG2;
  output N1BEG3;
  output N2BEG0;
  output N2BEG1;
  output N2BEG2;
  output N2BEG3;
  output N2BEG4;
  output N2BEG5;
  output N2BEG6;
  output N2BEG7;
  output N2BEGb0;
  output N2BEGb1;
  output N2BEGb2;
  output N2BEGb3;
  output N2BEGb4;
  output N2BEGb5;
  output N2BEGb6;
  output N2BEGb7;
  output N4BEG0;
  output N4BEG1;
  output N4BEG2;
  output N4BEG3;
  output NN4BEG0;
  output NN4BEG1;
  output NN4BEG2;
  output NN4BEG3;
  output E1BEG0;
  output E1BEG1;
  output E1BEG2;
  output E1BEG3;
  output E2BEG0;
  output E2BEG1;
  output E2BEG2;
  output E2BEG3;
  output E2BEG4;
  output E2BEG5;
  output E2BEG6;
  output E2BEG7;
  output E2BEGb0;
  output E2BEGb1;
  output E2BEGb2;
  output E2BEGb3;
  output E2BEGb4;
  output E2BEGb5;
  output E2BEGb6;
  output E2BEGb7;
  output EE4BEG0;
  output EE4BEG1;
  output EE4BEG2;
  output EE4BEG3;
  output E6BEG0;
  output E6BEG1;
  output S1BEG0;
  output S1BEG1;
  output S1BEG2;
  output S1BEG3;
  output S2BEG0;
  output S2BEG1;
  output S2BEG2;
  output S2BEG3;
  output S2BEG4;
  output S2BEG5;
  output S2BEG6;
  output S2BEG7;
  output S2BEGb0;
  output S2BEGb1;
  output S2BEGb2;
  output S2BEGb3;
  output S2BEGb4;
  output S2BEGb5;
  output S2BEGb6;
  output S2BEGb7;
  output S4BEG0;
  output S4BEG1;
  output S4BEG2;
  output S4BEG3;
  output SS4BEG0;
  output SS4BEG1;
  output SS4BEG2;
  output SS4BEG3;
  output W1BEG0;
  output W1BEG1;
  output W1BEG2;
  output W1BEG3;
  output W2BEG0;
  output W2BEG1;
  output W2BEG2;
  output W2BEG3;
  output W2BEG4;
  output W2BEG5;
  output W2BEG6;
  output W2BEG7;
  output W2BEGb0;
  output W2BEGb1;
  output W2BEGb2;
  output W2BEGb3;
  output W2BEGb4;
  output W2BEGb5;
  output W2BEGb6;
  output W2BEGb7;
  output WW4BEG0;
  output WW4BEG1;
  output WW4BEG2;
  output WW4BEG3;
  output W6BEG0;
  output W6BEG1;
  output D0;
  output D1;
  output D2;
  output D3;
  output W_ADR0;
  output W_ADR1;
  output W_ADR2;
  output W_ADR3;
  output W_ADR4;
  output W_en;
  output A_ADR0;
  output A_ADR1;
  output A_ADR2;
  output A_ADR3;
  output A_ADR4;
  output B_ADR0;
  output B_ADR1;
  output B_ADR2;
  output B_ADR3;
  output B_ADR4;
  output J2MID_ABa_BEG0;
  output J2MID_ABa_BEG1;
  output J2MID_ABa_BEG2;
  output J2MID_ABa_BEG3;
  output J2MID_CDa_BEG0;
  output J2MID_CDa_BEG1;
  output J2MID_CDa_BEG2;
  output J2MID_CDa_BEG3;
  output J2MID_EFa_BEG0;
  output J2MID_EFa_BEG1;
  output J2MID_EFa_BEG2;
  output J2MID_EFa_BEG3;
  output J2MID_GHa_BEG0;
  output J2MID_GHa_BEG1;
  output J2MID_GHa_BEG2;
  output J2MID_GHa_BEG3;
  output J2MID_ABb_BEG0;
  output J2MID_ABb_BEG1;
  output J2MID_ABb_BEG2;
  output J2MID_ABb_BEG3;
  output J2MID_CDb_BEG0;
  output J2MID_CDb_BEG1;
  output J2MID_CDb_BEG2;
  output J2MID_CDb_BEG3;
  output J2MID_EFb_BEG0;
  output J2MID_EFb_BEG1;
  output J2MID_EFb_BEG2;
  output J2MID_EFb_BEG3;
  output J2MID_GHb_BEG0;
  output J2MID_GHb_BEG1;
  output J2MID_GHb_BEG2;
  output J2MID_GHb_BEG3;
  output J2END_AB_BEG0;
  output J2END_AB_BEG1;
  output J2END_AB_BEG2;
  output J2END_AB_BEG3;
  output J2END_CD_BEG0;
  output J2END_CD_BEG1;
  output J2END_CD_BEG2;
  output J2END_CD_BEG3;
  output J2END_EF_BEG0;
  output J2END_EF_BEG1;
  output J2END_EF_BEG2;
  output J2END_EF_BEG3;
  output J2END_GH_BEG0;
  output J2END_GH_BEG1;
  output J2END_GH_BEG2;
  output J2END_GH_BEG3;
  output JN2BEG0;
  output JN2BEG1;
  output JN2BEG2;
  output JN2BEG3;
  output JN2BEG4;
  output JN2BEG5;
  output JN2BEG6;
  output JN2BEG7;
  output JE2BEG0;
  output JE2BEG1;
  output JE2BEG2;
  output JE2BEG3;
  output JE2BEG4;
  output JE2BEG5;
  output JE2BEG6;
  output JE2BEG7;
  output JS2BEG0;
  output JS2BEG1;
  output JS2BEG2;
  output JS2BEG3;
  output JS2BEG4;
  output JS2BEG5;
  output JS2BEG6;
  output JS2BEG7;
  output JW2BEG0;
  output JW2BEG1;
  output JW2BEG2;
  output JW2BEG3;
  output JW2BEG4;
  output JW2BEG5;
  output JW2BEG6;
  output JW2BEG7;
  output J_l_AB_BEG0;
  output J_l_AB_BEG1;
  output J_l_AB_BEG2;
  output J_l_AB_BEG3;
  output J_l_CD_BEG0;
  output J_l_CD_BEG1;
  output J_l_CD_BEG2;
  output J_l_CD_BEG3;
  output J_l_EF_BEG0;
  output J_l_EF_BEG1;
  output J_l_EF_BEG2;
  output J_l_EF_BEG3;
  output J_l_GH_BEG0;
  output J_l_GH_BEG1;
  output J_l_GH_BEG2;
  output J_l_GH_BEG3;
  //global
  input [NoConfigBits-1:0] ConfigBits;
  input [NoConfigBits-1:0] ConfigBits_N;

  parameter GND0 = 1'b0;
  parameter GND = 1'b0;
  parameter VCC0 = 1'b1;
  parameter VCC = 1'b1;
  parameter VDD0 = 1'b1;
  parameter VDD = 1'b1;

  wire [ 4-1:0] N1BEG0_input;
  wire [ 4-1:0] N1BEG1_input;
  wire [ 4-1:0] N1BEG2_input;
  wire [ 4-1:0] N1BEG3_input;
  wire [ 1-1:0] N2BEG0_input;
  wire [ 1-1:0] N2BEG1_input;
  wire [ 1-1:0] N2BEG2_input;
  wire [ 1-1:0] N2BEG3_input;
  wire [ 1-1:0] N2BEG4_input;
  wire [ 1-1:0] N2BEG5_input;
  wire [ 1-1:0] N2BEG6_input;
  wire [ 1-1:0] N2BEG7_input;
  wire [ 1-1:0] N2BEGb0_input;
  wire [ 1-1:0] N2BEGb1_input;
  wire [ 1-1:0] N2BEGb2_input;
  wire [ 1-1:0] N2BEGb3_input;
  wire [ 1-1:0] N2BEGb4_input;
  wire [ 1-1:0] N2BEGb5_input;
  wire [ 1-1:0] N2BEGb6_input;
  wire [ 1-1:0] N2BEGb7_input;
  wire [ 4-1:0] N4BEG0_input;
  wire [ 4-1:0] N4BEG1_input;
  wire [ 4-1:0] N4BEG2_input;
  wire [ 4-1:0] N4BEG3_input;
  wire [ 8-1:0] NN4BEG0_input;
  wire [ 8-1:0] NN4BEG1_input;
  wire [ 8-1:0] NN4BEG2_input;
  wire [ 8-1:0] NN4BEG3_input;
  wire [ 4-1:0] E1BEG0_input;
  wire [ 4-1:0] E1BEG1_input;
  wire [ 4-1:0] E1BEG2_input;
  wire [ 4-1:0] E1BEG3_input;
  wire [ 1-1:0] E2BEG0_input;
  wire [ 1-1:0] E2BEG1_input;
  wire [ 1-1:0] E2BEG2_input;
  wire [ 1-1:0] E2BEG3_input;
  wire [ 1-1:0] E2BEG4_input;
  wire [ 1-1:0] E2BEG5_input;
  wire [ 1-1:0] E2BEG6_input;
  wire [ 1-1:0] E2BEG7_input;
  wire [ 1-1:0] E2BEGb0_input;
  wire [ 1-1:0] E2BEGb1_input;
  wire [ 1-1:0] E2BEGb2_input;
  wire [ 1-1:0] E2BEGb3_input;
  wire [ 1-1:0] E2BEGb4_input;
  wire [ 1-1:0] E2BEGb5_input;
  wire [ 1-1:0] E2BEGb6_input;
  wire [ 1-1:0] E2BEGb7_input;
  wire [ 8-1:0] EE4BEG0_input;
  wire [ 8-1:0] EE4BEG1_input;
  wire [ 8-1:0] EE4BEG2_input;
  wire [ 8-1:0] EE4BEG3_input;
  wire [16-1:0] E6BEG0_input;
  wire [16-1:0] E6BEG1_input;
  wire [ 4-1:0] S1BEG0_input;
  wire [ 4-1:0] S1BEG1_input;
  wire [ 4-1:0] S1BEG2_input;
  wire [ 4-1:0] S1BEG3_input;
  wire [ 1-1:0] S2BEG0_input;
  wire [ 1-1:0] S2BEG1_input;
  wire [ 1-1:0] S2BEG2_input;
  wire [ 1-1:0] S2BEG3_input;
  wire [ 1-1:0] S2BEG4_input;
  wire [ 1-1:0] S2BEG5_input;
  wire [ 1-1:0] S2BEG6_input;
  wire [ 1-1:0] S2BEG7_input;
  wire [ 1-1:0] S2BEGb0_input;
  wire [ 1-1:0] S2BEGb1_input;
  wire [ 1-1:0] S2BEGb2_input;
  wire [ 1-1:0] S2BEGb3_input;
  wire [ 1-1:0] S2BEGb4_input;
  wire [ 1-1:0] S2BEGb5_input;
  wire [ 1-1:0] S2BEGb6_input;
  wire [ 1-1:0] S2BEGb7_input;
  wire [ 4-1:0] S4BEG0_input;
  wire [ 4-1:0] S4BEG1_input;
  wire [ 4-1:0] S4BEG2_input;
  wire [ 4-1:0] S4BEG3_input;
  wire [ 8-1:0] SS4BEG0_input;
  wire [ 8-1:0] SS4BEG1_input;
  wire [ 8-1:0] SS4BEG2_input;
  wire [ 8-1:0] SS4BEG3_input;
  wire [ 4-1:0] W1BEG0_input;
  wire [ 4-1:0] W1BEG1_input;
  wire [ 4-1:0] W1BEG2_input;
  wire [ 4-1:0] W1BEG3_input;
  wire [ 1-1:0] W2BEG0_input;
  wire [ 1-1:0] W2BEG1_input;
  wire [ 1-1:0] W2BEG2_input;
  wire [ 1-1:0] W2BEG3_input;
  wire [ 1-1:0] W2BEG4_input;
  wire [ 1-1:0] W2BEG5_input;
  wire [ 1-1:0] W2BEG6_input;
  wire [ 1-1:0] W2BEG7_input;
  wire [ 1-1:0] W2BEGb0_input;
  wire [ 1-1:0] W2BEGb1_input;
  wire [ 1-1:0] W2BEGb2_input;
  wire [ 1-1:0] W2BEGb3_input;
  wire [ 1-1:0] W2BEGb4_input;
  wire [ 1-1:0] W2BEGb5_input;
  wire [ 1-1:0] W2BEGb6_input;
  wire [ 1-1:0] W2BEGb7_input;
  wire [ 8-1:0] WW4BEG0_input;
  wire [ 8-1:0] WW4BEG1_input;
  wire [ 8-1:0] WW4BEG2_input;
  wire [ 8-1:0] WW4BEG3_input;
  wire [16-1:0] W6BEG0_input;
  wire [16-1:0] W6BEG1_input;
  wire [ 4-1:0] D0_input;
  wire [ 4-1:0] D1_input;
  wire [ 4-1:0] D2_input;
  wire [ 4-1:0] D3_input;
  wire [ 4-1:0] W_ADR0_input;
  wire [ 4-1:0] W_ADR1_input;
  wire [ 4-1:0] W_ADR2_input;
  wire [ 4-1:0] W_ADR3_input;
  wire [ 8-1:0] W_ADR4_input;
  wire [ 8-1:0] W_en_input;
  wire [ 4-1:0] A_ADR0_input;
  wire [ 4-1:0] A_ADR1_input;
  wire [ 4-1:0] A_ADR2_input;
  wire [ 4-1:0] A_ADR3_input;
  wire [ 8-1:0] A_ADR4_input;
  wire [ 4-1:0] B_ADR0_input;
  wire [ 4-1:0] B_ADR1_input;
  wire [ 4-1:0] B_ADR2_input;
  wire [ 4-1:0] B_ADR3_input;
  wire [ 8-1:0] B_ADR4_input;
  wire [ 4-1:0] J2MID_ABa_BEG0_input;
  wire [ 4-1:0] J2MID_ABa_BEG1_input;
  wire [ 4-1:0] J2MID_ABa_BEG2_input;
  wire [ 4-1:0] J2MID_ABa_BEG3_input;
  wire [ 4-1:0] J2MID_CDa_BEG0_input;
  wire [ 4-1:0] J2MID_CDa_BEG1_input;
  wire [ 4-1:0] J2MID_CDa_BEG2_input;
  wire [ 4-1:0] J2MID_CDa_BEG3_input;
  wire [ 4-1:0] J2MID_EFa_BEG0_input;
  wire [ 4-1:0] J2MID_EFa_BEG1_input;
  wire [ 4-1:0] J2MID_EFa_BEG2_input;
  wire [ 4-1:0] J2MID_EFa_BEG3_input;
  wire [ 4-1:0] J2MID_GHa_BEG0_input;
  wire [ 4-1:0] J2MID_GHa_BEG1_input;
  wire [ 4-1:0] J2MID_GHa_BEG2_input;
  wire [ 4-1:0] J2MID_GHa_BEG3_input;
  wire [ 4-1:0] J2MID_ABb_BEG0_input;
  wire [ 4-1:0] J2MID_ABb_BEG1_input;
  wire [ 4-1:0] J2MID_ABb_BEG2_input;
  wire [ 4-1:0] J2MID_ABb_BEG3_input;
  wire [ 4-1:0] J2MID_CDb_BEG0_input;
  wire [ 4-1:0] J2MID_CDb_BEG1_input;
  wire [ 4-1:0] J2MID_CDb_BEG2_input;
  wire [ 4-1:0] J2MID_CDb_BEG3_input;
  wire [ 4-1:0] J2MID_EFb_BEG0_input;
  wire [ 4-1:0] J2MID_EFb_BEG1_input;
  wire [ 4-1:0] J2MID_EFb_BEG2_input;
  wire [ 4-1:0] J2MID_EFb_BEG3_input;
  wire [ 4-1:0] J2MID_GHb_BEG0_input;
  wire [ 4-1:0] J2MID_GHb_BEG1_input;
  wire [ 4-1:0] J2MID_GHb_BEG2_input;
  wire [ 4-1:0] J2MID_GHb_BEG3_input;
  wire [ 4-1:0] J2END_AB_BEG0_input;
  wire [ 4-1:0] J2END_AB_BEG1_input;
  wire [ 4-1:0] J2END_AB_BEG2_input;
  wire [ 4-1:0] J2END_AB_BEG3_input;
  wire [ 4-1:0] J2END_CD_BEG0_input;
  wire [ 4-1:0] J2END_CD_BEG1_input;
  wire [ 4-1:0] J2END_CD_BEG2_input;
  wire [ 4-1:0] J2END_CD_BEG3_input;
  wire [ 4-1:0] J2END_EF_BEG0_input;
  wire [ 4-1:0] J2END_EF_BEG1_input;
  wire [ 4-1:0] J2END_EF_BEG2_input;
  wire [ 4-1:0] J2END_EF_BEG3_input;
  wire [ 4-1:0] J2END_GH_BEG0_input;
  wire [ 4-1:0] J2END_GH_BEG1_input;
  wire [ 4-1:0] J2END_GH_BEG2_input;
  wire [ 4-1:0] J2END_GH_BEG3_input;
  wire [16-1:0] JN2BEG0_input;
  wire [16-1:0] JN2BEG1_input;
  wire [16-1:0] JN2BEG2_input;
  wire [16-1:0] JN2BEG3_input;
  wire [16-1:0] JN2BEG4_input;
  wire [16-1:0] JN2BEG5_input;
  wire [16-1:0] JN2BEG6_input;
  wire [16-1:0] JN2BEG7_input;
  wire [16-1:0] JE2BEG0_input;
  wire [16-1:0] JE2BEG1_input;
  wire [16-1:0] JE2BEG2_input;
  wire [16-1:0] JE2BEG3_input;
  wire [16-1:0] JE2BEG4_input;
  wire [16-1:0] JE2BEG5_input;
  wire [16-1:0] JE2BEG6_input;
  wire [16-1:0] JE2BEG7_input;
  wire [16-1:0] JS2BEG0_input;
  wire [16-1:0] JS2BEG1_input;
  wire [16-1:0] JS2BEG2_input;
  wire [16-1:0] JS2BEG3_input;
  wire [16-1:0] JS2BEG4_input;
  wire [16-1:0] JS2BEG5_input;
  wire [16-1:0] JS2BEG6_input;
  wire [16-1:0] JS2BEG7_input;
  wire [16-1:0] JW2BEG0_input;
  wire [16-1:0] JW2BEG1_input;
  wire [16-1:0] JW2BEG2_input;
  wire [16-1:0] JW2BEG3_input;
  wire [16-1:0] JW2BEG4_input;
  wire [16-1:0] JW2BEG5_input;
  wire [16-1:0] JW2BEG6_input;
  wire [16-1:0] JW2BEG7_input;
  wire [ 4-1:0] J_l_AB_BEG0_input;
  wire [ 4-1:0] J_l_AB_BEG1_input;
  wire [ 4-1:0] J_l_AB_BEG2_input;
  wire [ 4-1:0] J_l_AB_BEG3_input;
  wire [ 4-1:0] J_l_CD_BEG0_input;
  wire [ 4-1:0] J_l_CD_BEG1_input;
  wire [ 4-1:0] J_l_CD_BEG2_input;
  wire [ 4-1:0] J_l_CD_BEG3_input;
  wire [ 4-1:0] J_l_EF_BEG0_input;
  wire [ 4-1:0] J_l_EF_BEG1_input;
  wire [ 4-1:0] J_l_EF_BEG2_input;
  wire [ 4-1:0] J_l_EF_BEG3_input;
  wire [ 4-1:0] J_l_GH_BEG0_input;
  wire [ 4-1:0] J_l_GH_BEG1_input;
  wire [ 4-1:0] J_l_GH_BEG2_input;
  wire [ 4-1:0] J_l_GH_BEG3_input;

  wire [ 2-1:0] DEBUG_select_N1BEG0;
  wire [ 2-1:0] DEBUG_select_N1BEG1;
  wire [ 2-1:0] DEBUG_select_N1BEG2;
  wire [ 2-1:0] DEBUG_select_N1BEG3;
  wire [ 2-1:0] DEBUG_select_N4BEG0;
  wire [ 2-1:0] DEBUG_select_N4BEG1;
  wire [ 2-1:0] DEBUG_select_N4BEG2;
  wire [ 2-1:0] DEBUG_select_N4BEG3;
  wire [ 3-1:0] DEBUG_select_NN4BEG0;
  wire [ 3-1:0] DEBUG_select_NN4BEG1;
  wire [ 3-1:0] DEBUG_select_NN4BEG2;
  wire [ 3-1:0] DEBUG_select_NN4BEG3;
  wire [ 2-1:0] DEBUG_select_E1BEG0;
  wire [ 2-1:0] DEBUG_select_E1BEG1;
  wire [ 2-1:0] DEBUG_select_E1BEG2;
  wire [ 2-1:0] DEBUG_select_E1BEG3;
  wire [ 3-1:0] DEBUG_select_EE4BEG0;
  wire [ 3-1:0] DEBUG_select_EE4BEG1;
  wire [ 3-1:0] DEBUG_select_EE4BEG2;
  wire [ 3-1:0] DEBUG_select_EE4BEG3;
  wire [ 4-1:0] DEBUG_select_E6BEG0;
  wire [ 4-1:0] DEBUG_select_E6BEG1;
  wire [ 2-1:0] DEBUG_select_S1BEG0;
  wire [ 2-1:0] DEBUG_select_S1BEG1;
  wire [ 2-1:0] DEBUG_select_S1BEG2;
  wire [ 2-1:0] DEBUG_select_S1BEG3;
  wire [ 2-1:0] DEBUG_select_S4BEG0;
  wire [ 2-1:0] DEBUG_select_S4BEG1;
  wire [ 2-1:0] DEBUG_select_S4BEG2;
  wire [ 2-1:0] DEBUG_select_S4BEG3;
  wire [ 3-1:0] DEBUG_select_SS4BEG0;
  wire [ 3-1:0] DEBUG_select_SS4BEG1;
  wire [ 3-1:0] DEBUG_select_SS4BEG2;
  wire [ 3-1:0] DEBUG_select_SS4BEG3;
  wire [ 2-1:0] DEBUG_select_W1BEG0;
  wire [ 2-1:0] DEBUG_select_W1BEG1;
  wire [ 2-1:0] DEBUG_select_W1BEG2;
  wire [ 2-1:0] DEBUG_select_W1BEG3;
  wire [ 3-1:0] DEBUG_select_WW4BEG0;
  wire [ 3-1:0] DEBUG_select_WW4BEG1;
  wire [ 3-1:0] DEBUG_select_WW4BEG2;
  wire [ 3-1:0] DEBUG_select_WW4BEG3;
  wire [ 4-1:0] DEBUG_select_W6BEG0;
  wire [ 4-1:0] DEBUG_select_W6BEG1;
  wire [ 2-1:0] DEBUG_select_D0;
  wire [ 2-1:0] DEBUG_select_D1;
  wire [ 2-1:0] DEBUG_select_D2;
  wire [ 2-1:0] DEBUG_select_D3;
  wire [ 2-1:0] DEBUG_select_W_ADR0;
  wire [ 2-1:0] DEBUG_select_W_ADR1;
  wire [ 2-1:0] DEBUG_select_W_ADR2;
  wire [ 2-1:0] DEBUG_select_W_ADR3;
  wire [ 3-1:0] DEBUG_select_W_ADR4;
  wire [ 3-1:0] DEBUG_select_W_en;
  wire [ 2-1:0] DEBUG_select_A_ADR0;
  wire [ 2-1:0] DEBUG_select_A_ADR1;
  wire [ 2-1:0] DEBUG_select_A_ADR2;
  wire [ 2-1:0] DEBUG_select_A_ADR3;
  wire [ 3-1:0] DEBUG_select_A_ADR4;
  wire [ 2-1:0] DEBUG_select_B_ADR0;
  wire [ 2-1:0] DEBUG_select_B_ADR1;
  wire [ 2-1:0] DEBUG_select_B_ADR2;
  wire [ 2-1:0] DEBUG_select_B_ADR3;
  wire [ 3-1:0] DEBUG_select_B_ADR4;
  wire [ 2-1:0] DEBUG_select_J2MID_ABa_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_ABa_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_ABa_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_ABa_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_CDa_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_CDa_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_CDa_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_CDa_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_EFa_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_EFa_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_EFa_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_EFa_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_GHa_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_GHa_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_GHa_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_GHa_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_ABb_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_ABb_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_ABb_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_ABb_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_CDb_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_CDb_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_CDb_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_CDb_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_EFb_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_EFb_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_EFb_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_EFb_BEG3;
  wire [ 2-1:0] DEBUG_select_J2MID_GHb_BEG0;
  wire [ 2-1:0] DEBUG_select_J2MID_GHb_BEG1;
  wire [ 2-1:0] DEBUG_select_J2MID_GHb_BEG2;
  wire [ 2-1:0] DEBUG_select_J2MID_GHb_BEG3;
  wire [ 2-1:0] DEBUG_select_J2END_AB_BEG0;
  wire [ 2-1:0] DEBUG_select_J2END_AB_BEG1;
  wire [ 2-1:0] DEBUG_select_J2END_AB_BEG2;
  wire [ 2-1:0] DEBUG_select_J2END_AB_BEG3;
  wire [ 2-1:0] DEBUG_select_J2END_CD_BEG0;
  wire [ 2-1:0] DEBUG_select_J2END_CD_BEG1;
  wire [ 2-1:0] DEBUG_select_J2END_CD_BEG2;
  wire [ 2-1:0] DEBUG_select_J2END_CD_BEG3;
  wire [ 2-1:0] DEBUG_select_J2END_EF_BEG0;
  wire [ 2-1:0] DEBUG_select_J2END_EF_BEG1;
  wire [ 2-1:0] DEBUG_select_J2END_EF_BEG2;
  wire [ 2-1:0] DEBUG_select_J2END_EF_BEG3;
  wire [ 2-1:0] DEBUG_select_J2END_GH_BEG0;
  wire [ 2-1:0] DEBUG_select_J2END_GH_BEG1;
  wire [ 2-1:0] DEBUG_select_J2END_GH_BEG2;
  wire [ 2-1:0] DEBUG_select_J2END_GH_BEG3;
  wire [ 4-1:0] DEBUG_select_JN2BEG0;
  wire [ 4-1:0] DEBUG_select_JN2BEG1;
  wire [ 4-1:0] DEBUG_select_JN2BEG2;
  wire [ 4-1:0] DEBUG_select_JN2BEG3;
  wire [ 4-1:0] DEBUG_select_JN2BEG4;
  wire [ 4-1:0] DEBUG_select_JN2BEG5;
  wire [ 4-1:0] DEBUG_select_JN2BEG6;
  wire [ 4-1:0] DEBUG_select_JN2BEG7;
  wire [ 4-1:0] DEBUG_select_JE2BEG0;
  wire [ 4-1:0] DEBUG_select_JE2BEG1;
  wire [ 4-1:0] DEBUG_select_JE2BEG2;
  wire [ 4-1:0] DEBUG_select_JE2BEG3;
  wire [ 4-1:0] DEBUG_select_JE2BEG4;
  wire [ 4-1:0] DEBUG_select_JE2BEG5;
  wire [ 4-1:0] DEBUG_select_JE2BEG6;
  wire [ 4-1:0] DEBUG_select_JE2BEG7;
  wire [ 4-1:0] DEBUG_select_JS2BEG0;
  wire [ 4-1:0] DEBUG_select_JS2BEG1;
  wire [ 4-1:0] DEBUG_select_JS2BEG2;
  wire [ 4-1:0] DEBUG_select_JS2BEG3;
  wire [ 4-1:0] DEBUG_select_JS2BEG4;
  wire [ 4-1:0] DEBUG_select_JS2BEG5;
  wire [ 4-1:0] DEBUG_select_JS2BEG6;
  wire [ 4-1:0] DEBUG_select_JS2BEG7;
  wire [ 4-1:0] DEBUG_select_JW2BEG0;
  wire [ 4-1:0] DEBUG_select_JW2BEG1;
  wire [ 4-1:0] DEBUG_select_JW2BEG2;
  wire [ 4-1:0] DEBUG_select_JW2BEG3;
  wire [ 4-1:0] DEBUG_select_JW2BEG4;
  wire [ 4-1:0] DEBUG_select_JW2BEG5;
  wire [ 4-1:0] DEBUG_select_JW2BEG6;
  wire [ 4-1:0] DEBUG_select_JW2BEG7;
  wire [ 2-1:0] DEBUG_select_J_l_AB_BEG0;
  wire [ 2-1:0] DEBUG_select_J_l_AB_BEG1;
  wire [ 2-1:0] DEBUG_select_J_l_AB_BEG2;
  wire [ 2-1:0] DEBUG_select_J_l_AB_BEG3;
  wire [ 2-1:0] DEBUG_select_J_l_CD_BEG0;
  wire [ 2-1:0] DEBUG_select_J_l_CD_BEG1;
  wire [ 2-1:0] DEBUG_select_J_l_CD_BEG2;
  wire [ 2-1:0] DEBUG_select_J_l_CD_BEG3;
  wire [ 2-1:0] DEBUG_select_J_l_EF_BEG0;
  wire [ 2-1:0] DEBUG_select_J_l_EF_BEG1;
  wire [ 2-1:0] DEBUG_select_J_l_EF_BEG2;
  wire [ 2-1:0] DEBUG_select_J_l_EF_BEG3;
  wire [ 2-1:0] DEBUG_select_J_l_GH_BEG0;
  wire [ 2-1:0] DEBUG_select_J_l_GH_BEG1;
  wire [ 2-1:0] DEBUG_select_J_l_GH_BEG2;
  wire [ 2-1:0] DEBUG_select_J_l_GH_BEG3;

  // The configuration bits (if any) are just a long shift register

  // This shift register is padded to an even number of flops/latches
  // switch matrix multiplexer  N1BEG0         MUX-4
  assign N1BEG0_input = {J_l_CD_END1, JW2END3, J2MID_CDb_END3, AD2};
  cus_mux41_buf inst_cus_mux41_buf_N1BEG0 (
      .A0 (N1BEG0_input[0]),
      .A1 (N1BEG0_input[1]),
      .A2 (N1BEG0_input[2]),
      .A3 (N1BEG0_input[3]),
      .S0 (ConfigBits[0+0]),
      .S0N(ConfigBits_N[0+0]),
      .S1 (ConfigBits[0+1]),
      .S1N(ConfigBits_N[0+1]),
      .X  (N1BEG0)
  );

  // switch matrix multiplexer  N1BEG1         MUX-4
  assign N1BEG1_input = {J_l_EF_END2, JW2END0, J2MID_EFb_END0, AD3};
  cus_mux41_buf inst_cus_mux41_buf_N1BEG1 (
      .A0 (N1BEG1_input[0]),
      .A1 (N1BEG1_input[1]),
      .A2 (N1BEG1_input[2]),
      .A3 (N1BEG1_input[3]),
      .S0 (ConfigBits[2+0]),
      .S0N(ConfigBits_N[2+0]),
      .S1 (ConfigBits[2+1]),
      .S1N(ConfigBits_N[2+1]),
      .X  (N1BEG1)
  );

  // switch matrix multiplexer  N1BEG2         MUX-4
  assign N1BEG2_input = {J_l_GH_END3, JW2END1, J2MID_GHb_END1, BD0};
  cus_mux41_buf inst_cus_mux41_buf_N1BEG2 (
      .A0 (N1BEG2_input[0]),
      .A1 (N1BEG2_input[1]),
      .A2 (N1BEG2_input[2]),
      .A3 (N1BEG2_input[3]),
      .S0 (ConfigBits[4+0]),
      .S0N(ConfigBits_N[4+0]),
      .S1 (ConfigBits[4+1]),
      .S1N(ConfigBits_N[4+1]),
      .X  (N1BEG2)
  );

  // switch matrix multiplexer  N1BEG3         MUX-4
  assign N1BEG3_input = {J_l_AB_END0, JW2END2, J2MID_ABb_END2, BD1};
  cus_mux41_buf inst_cus_mux41_buf_N1BEG3 (
      .A0 (N1BEG3_input[0]),
      .A1 (N1BEG3_input[1]),
      .A2 (N1BEG3_input[2]),
      .A3 (N1BEG3_input[3]),
      .S0 (ConfigBits[6+0]),
      .S0N(ConfigBits_N[6+0]),
      .S1 (ConfigBits[6+1]),
      .S1N(ConfigBits_N[6+1]),
      .X  (N1BEG3)
  );

  // switch matrix multiplexer  N2BEG0         MUX-1
  assign N2BEG0 = JN2END0;
  // switch matrix multiplexer  N2BEG1         MUX-1
  assign N2BEG1 = JN2END1;
  // switch matrix multiplexer  N2BEG2         MUX-1
  assign N2BEG2 = JN2END2;
  // switch matrix multiplexer  N2BEG3         MUX-1
  assign N2BEG3 = JN2END3;
  // switch matrix multiplexer  N2BEG4         MUX-1
  assign N2BEG4 = JN2END4;
  // switch matrix multiplexer  N2BEG5         MUX-1
  assign N2BEG5 = JN2END5;
  // switch matrix multiplexer  N2BEG6         MUX-1
  assign N2BEG6 = JN2END6;
  // switch matrix multiplexer  N2BEG7         MUX-1
  assign N2BEG7 = JN2END7;
  // switch matrix multiplexer  N2BEGb0         MUX-1
  assign N2BEGb0 = N2MID0;
  // switch matrix multiplexer  N2BEGb1         MUX-1
  assign N2BEGb1 = N2MID1;
  // switch matrix multiplexer  N2BEGb2         MUX-1
  assign N2BEGb2 = N2MID2;
  // switch matrix multiplexer  N2BEGb3         MUX-1
  assign N2BEGb3 = N2MID3;
  // switch matrix multiplexer  N2BEGb4         MUX-1
  assign N2BEGb4 = N2MID4;
  // switch matrix multiplexer  N2BEGb5         MUX-1
  assign N2BEGb5 = N2MID5;
  // switch matrix multiplexer  N2BEGb6         MUX-1
  assign N2BEGb6 = N2MID6;
  // switch matrix multiplexer  N2BEGb7         MUX-1
  assign N2BEGb7 = N2MID7;
  // switch matrix multiplexer  N4BEG0         MUX-4
  assign N4BEG0_input = {BD0, E6END1, N4END1, N2END2};
  cus_mux41_buf inst_cus_mux41_buf_N4BEG0 (
      .A0 (N4BEG0_input[0]),
      .A1 (N4BEG0_input[1]),
      .A2 (N4BEG0_input[2]),
      .A3 (N4BEG0_input[3]),
      .S0 (ConfigBits[8+0]),
      .S0N(ConfigBits_N[8+0]),
      .S1 (ConfigBits[8+1]),
      .S1N(ConfigBits_N[8+1]),
      .X  (N4BEG0)
  );

  // switch matrix multiplexer  N4BEG1         MUX-4
  assign N4BEG1_input = {BD1, E6END0, N4END2, N2END3};
  cus_mux41_buf inst_cus_mux41_buf_N4BEG1 (
      .A0 (N4BEG1_input[0]),
      .A1 (N4BEG1_input[1]),
      .A2 (N4BEG1_input[2]),
      .A3 (N4BEG1_input[3]),
      .S0 (ConfigBits[10+0]),
      .S0N(ConfigBits_N[10+0]),
      .S1 (ConfigBits[10+1]),
      .S1N(ConfigBits_N[10+1]),
      .X  (N4BEG1)
  );

  // switch matrix multiplexer  N4BEG2         MUX-4
  assign N4BEG2_input = {BD2, W6END1, N4END3, N2END0};
  cus_mux41_buf inst_cus_mux41_buf_N4BEG2 (
      .A0 (N4BEG2_input[0]),
      .A1 (N4BEG2_input[1]),
      .A2 (N4BEG2_input[2]),
      .A3 (N4BEG2_input[3]),
      .S0 (ConfigBits[12+0]),
      .S0N(ConfigBits_N[12+0]),
      .S1 (ConfigBits[12+1]),
      .S1N(ConfigBits_N[12+1]),
      .X  (N4BEG2)
  );

  // switch matrix multiplexer  N4BEG3         MUX-4
  assign N4BEG3_input = {BD3, W6END0, N4END0, N2END1};
  cus_mux41_buf inst_cus_mux41_buf_N4BEG3 (
      .A0 (N4BEG3_input[0]),
      .A1 (N4BEG3_input[1]),
      .A2 (N4BEG3_input[2]),
      .A3 (N4BEG3_input[3]),
      .S0 (ConfigBits[14+0]),
      .S0N(ConfigBits_N[14+0]),
      .S1 (ConfigBits[14+1]),
      .S1N(ConfigBits_N[14+1]),
      .X  (N4BEG3)
  );

  // switch matrix multiplexer  NN4BEG0         MUX-8
  assign NN4BEG0_input = {
    J2END_GH_END1, J2MID_CDb_END1, J2MID_ABb_END1, BD1, AD1, W1END2, E1END2, N1END2
  };
  cus_mux81_buf inst_cus_mux81_buf_NN4BEG0 (
      .A0 (NN4BEG0_input[0]),
      .A1 (NN4BEG0_input[1]),
      .A2 (NN4BEG0_input[2]),
      .A3 (NN4BEG0_input[3]),
      .A4 (NN4BEG0_input[4]),
      .A5 (NN4BEG0_input[5]),
      .A6 (NN4BEG0_input[6]),
      .A7 (NN4BEG0_input[7]),
      .S0 (ConfigBits[16+0]),
      .S0N(ConfigBits_N[16+0]),
      .S1 (ConfigBits[16+1]),
      .S1N(ConfigBits_N[16+1]),
      .S2 (ConfigBits[16+2]),
      .S2N(ConfigBits_N[16+2]),
      .X  (NN4BEG0)
  );

  // switch matrix multiplexer  NN4BEG1         MUX-8
  assign NN4BEG1_input = {
    J2END_EF_END1, J2MID_CDa_END2, J2MID_ABa_END2, BD2, AD2, W1END3, E1END3, N1END3
  };
  cus_mux81_buf inst_cus_mux81_buf_NN4BEG1 (
      .A0 (NN4BEG1_input[0]),
      .A1 (NN4BEG1_input[1]),
      .A2 (NN4BEG1_input[2]),
      .A3 (NN4BEG1_input[3]),
      .A4 (NN4BEG1_input[4]),
      .A5 (NN4BEG1_input[5]),
      .A6 (NN4BEG1_input[6]),
      .A7 (NN4BEG1_input[7]),
      .S0 (ConfigBits[19+0]),
      .S0N(ConfigBits_N[19+0]),
      .S1 (ConfigBits[19+1]),
      .S1N(ConfigBits_N[19+1]),
      .S2 (ConfigBits[19+2]),
      .S2N(ConfigBits_N[19+2]),
      .X  (NN4BEG1)
  );

  // switch matrix multiplexer  NN4BEG2         MUX-8
  assign NN4BEG2_input = {
    J2END_CD_END1, J2MID_GHb_END1, J2MID_EFb_END1, BD3, AD3, W1END0, E1END0, N1END0
  };
  cus_mux81_buf inst_cus_mux81_buf_NN4BEG2 (
      .A0 (NN4BEG2_input[0]),
      .A1 (NN4BEG2_input[1]),
      .A2 (NN4BEG2_input[2]),
      .A3 (NN4BEG2_input[3]),
      .A4 (NN4BEG2_input[4]),
      .A5 (NN4BEG2_input[5]),
      .A6 (NN4BEG2_input[6]),
      .A7 (NN4BEG2_input[7]),
      .S0 (ConfigBits[22+0]),
      .S0N(ConfigBits_N[22+0]),
      .S1 (ConfigBits[22+1]),
      .S1N(ConfigBits_N[22+1]),
      .S2 (ConfigBits[22+2]),
      .S2N(ConfigBits_N[22+2]),
      .X  (NN4BEG2)
  );

  // switch matrix multiplexer  NN4BEG3         MUX-8
  assign NN4BEG3_input = {
    J2END_AB_END1, J2MID_GHa_END2, J2MID_EFa_END2, BD0, AD0, W1END1, E1END1, N1END1
  };
  cus_mux81_buf inst_cus_mux81_buf_NN4BEG3 (
      .A0 (NN4BEG3_input[0]),
      .A1 (NN4BEG3_input[1]),
      .A2 (NN4BEG3_input[2]),
      .A3 (NN4BEG3_input[3]),
      .A4 (NN4BEG3_input[4]),
      .A5 (NN4BEG3_input[5]),
      .A6 (NN4BEG3_input[6]),
      .A7 (NN4BEG3_input[7]),
      .S0 (ConfigBits[25+0]),
      .S0N(ConfigBits_N[25+0]),
      .S1 (ConfigBits[25+1]),
      .S1N(ConfigBits_N[25+1]),
      .S2 (ConfigBits[25+2]),
      .S2N(ConfigBits_N[25+2]),
      .X  (NN4BEG3)
  );

  // switch matrix multiplexer  E1BEG0         MUX-4
  assign E1BEG0_input = {J_l_CD_END1, JN2END3, J2MID_CDb_END3, AD3};
  cus_mux41_buf inst_cus_mux41_buf_E1BEG0 (
      .A0 (E1BEG0_input[0]),
      .A1 (E1BEG0_input[1]),
      .A2 (E1BEG0_input[2]),
      .A3 (E1BEG0_input[3]),
      .S0 (ConfigBits[28+0]),
      .S0N(ConfigBits_N[28+0]),
      .S1 (ConfigBits[28+1]),
      .S1N(ConfigBits_N[28+1]),
      .X  (E1BEG0)
  );

  // switch matrix multiplexer  E1BEG1         MUX-4
  assign E1BEG1_input = {J_l_EF_END2, JN2END0, J2MID_EFb_END0, BD0};
  cus_mux41_buf inst_cus_mux41_buf_E1BEG1 (
      .A0 (E1BEG1_input[0]),
      .A1 (E1BEG1_input[1]),
      .A2 (E1BEG1_input[2]),
      .A3 (E1BEG1_input[3]),
      .S0 (ConfigBits[30+0]),
      .S0N(ConfigBits_N[30+0]),
      .S1 (ConfigBits[30+1]),
      .S1N(ConfigBits_N[30+1]),
      .X  (E1BEG1)
  );

  // switch matrix multiplexer  E1BEG2         MUX-4
  assign E1BEG2_input = {J_l_GH_END3, JN2END1, J2MID_GHb_END1, BD1};
  cus_mux41_buf inst_cus_mux41_buf_E1BEG2 (
      .A0 (E1BEG2_input[0]),
      .A1 (E1BEG2_input[1]),
      .A2 (E1BEG2_input[2]),
      .A3 (E1BEG2_input[3]),
      .S0 (ConfigBits[32+0]),
      .S0N(ConfigBits_N[32+0]),
      .S1 (ConfigBits[32+1]),
      .S1N(ConfigBits_N[32+1]),
      .X  (E1BEG2)
  );

  // switch matrix multiplexer  E1BEG3         MUX-4
  assign E1BEG3_input = {J_l_AB_END0, JN2END2, J2MID_ABb_END2, BD2};
  cus_mux41_buf inst_cus_mux41_buf_E1BEG3 (
      .A0 (E1BEG3_input[0]),
      .A1 (E1BEG3_input[1]),
      .A2 (E1BEG3_input[2]),
      .A3 (E1BEG3_input[3]),
      .S0 (ConfigBits[34+0]),
      .S0N(ConfigBits_N[34+0]),
      .S1 (ConfigBits[34+1]),
      .S1N(ConfigBits_N[34+1]),
      .X  (E1BEG3)
  );

  // switch matrix multiplexer  E2BEG0         MUX-1
  assign E2BEG0 = JE2END0;
  // switch matrix multiplexer  E2BEG1         MUX-1
  assign E2BEG1 = JE2END1;
  // switch matrix multiplexer  E2BEG2         MUX-1
  assign E2BEG2 = JE2END2;
  // switch matrix multiplexer  E2BEG3         MUX-1
  assign E2BEG3 = JE2END3;
  // switch matrix multiplexer  E2BEG4         MUX-1
  assign E2BEG4 = JE2END4;
  // switch matrix multiplexer  E2BEG5         MUX-1
  assign E2BEG5 = JE2END5;
  // switch matrix multiplexer  E2BEG6         MUX-1
  assign E2BEG6 = JE2END6;
  // switch matrix multiplexer  E2BEG7         MUX-1
  assign E2BEG7 = JE2END7;
  // switch matrix multiplexer  E2BEGb0         MUX-1
  assign E2BEGb0 = E2MID0;
  // switch matrix multiplexer  E2BEGb1         MUX-1
  assign E2BEGb1 = E2MID1;
  // switch matrix multiplexer  E2BEGb2         MUX-1
  assign E2BEGb2 = E2MID2;
  // switch matrix multiplexer  E2BEGb3         MUX-1
  assign E2BEGb3 = E2MID3;
  // switch matrix multiplexer  E2BEGb4         MUX-1
  assign E2BEGb4 = E2MID4;
  // switch matrix multiplexer  E2BEGb5         MUX-1
  assign E2BEGb5 = E2MID5;
  // switch matrix multiplexer  E2BEGb6         MUX-1
  assign E2BEGb6 = E2MID6;
  // switch matrix multiplexer  E2BEGb7         MUX-1
  assign E2BEGb7 = E2MID7;
  // switch matrix multiplexer  EE4BEG0         MUX-8
  assign EE4BEG0_input = {
    J2END_GH_END0, J2MID_CDb_END1, J2MID_ABb_END1, BD1, AD1, S1END2, E1END2, N1END2
  };
  cus_mux81_buf inst_cus_mux81_buf_EE4BEG0 (
      .A0 (EE4BEG0_input[0]),
      .A1 (EE4BEG0_input[1]),
      .A2 (EE4BEG0_input[2]),
      .A3 (EE4BEG0_input[3]),
      .A4 (EE4BEG0_input[4]),
      .A5 (EE4BEG0_input[5]),
      .A6 (EE4BEG0_input[6]),
      .A7 (EE4BEG0_input[7]),
      .S0 (ConfigBits[36+0]),
      .S0N(ConfigBits_N[36+0]),
      .S1 (ConfigBits[36+1]),
      .S1N(ConfigBits_N[36+1]),
      .S2 (ConfigBits[36+2]),
      .S2N(ConfigBits_N[36+2]),
      .X  (EE4BEG0)
  );

  // switch matrix multiplexer  EE4BEG1         MUX-8
  assign EE4BEG1_input = {
    J2END_EF_END0, J2MID_CDa_END2, J2MID_ABa_END2, BD2, AD2, S1END3, E1END3, N1END3
  };
  cus_mux81_buf inst_cus_mux81_buf_EE4BEG1 (
      .A0 (EE4BEG1_input[0]),
      .A1 (EE4BEG1_input[1]),
      .A2 (EE4BEG1_input[2]),
      .A3 (EE4BEG1_input[3]),
      .A4 (EE4BEG1_input[4]),
      .A5 (EE4BEG1_input[5]),
      .A6 (EE4BEG1_input[6]),
      .A7 (EE4BEG1_input[7]),
      .S0 (ConfigBits[39+0]),
      .S0N(ConfigBits_N[39+0]),
      .S1 (ConfigBits[39+1]),
      .S1N(ConfigBits_N[39+1]),
      .S2 (ConfigBits[39+2]),
      .S2N(ConfigBits_N[39+2]),
      .X  (EE4BEG1)
  );

  // switch matrix multiplexer  EE4BEG2         MUX-8
  assign EE4BEG2_input = {
    J2END_CD_END0, J2MID_GHb_END1, J2MID_EFb_END1, BD3, AD3, S1END0, E1END0, N1END0
  };
  cus_mux81_buf inst_cus_mux81_buf_EE4BEG2 (
      .A0 (EE4BEG2_input[0]),
      .A1 (EE4BEG2_input[1]),
      .A2 (EE4BEG2_input[2]),
      .A3 (EE4BEG2_input[3]),
      .A4 (EE4BEG2_input[4]),
      .A5 (EE4BEG2_input[5]),
      .A6 (EE4BEG2_input[6]),
      .A7 (EE4BEG2_input[7]),
      .S0 (ConfigBits[42+0]),
      .S0N(ConfigBits_N[42+0]),
      .S1 (ConfigBits[42+1]),
      .S1N(ConfigBits_N[42+1]),
      .S2 (ConfigBits[42+2]),
      .S2N(ConfigBits_N[42+2]),
      .X  (EE4BEG2)
  );

  // switch matrix multiplexer  EE4BEG3         MUX-8
  assign EE4BEG3_input = {
    J2END_AB_END0, J2MID_GHa_END2, J2MID_EFa_END2, BD0, AD0, S1END1, E1END1, N1END1
  };
  cus_mux81_buf inst_cus_mux81_buf_EE4BEG3 (
      .A0 (EE4BEG3_input[0]),
      .A1 (EE4BEG3_input[1]),
      .A2 (EE4BEG3_input[2]),
      .A3 (EE4BEG3_input[3]),
      .A4 (EE4BEG3_input[4]),
      .A5 (EE4BEG3_input[5]),
      .A6 (EE4BEG3_input[6]),
      .A7 (EE4BEG3_input[7]),
      .S0 (ConfigBits[45+0]),
      .S0N(ConfigBits_N[45+0]),
      .S1 (ConfigBits[45+1]),
      .S1N(ConfigBits_N[45+1]),
      .S2 (ConfigBits[45+2]),
      .S2N(ConfigBits_N[45+2]),
      .X  (EE4BEG3)
  );

  // switch matrix multiplexer  E6BEG0         MUX-16
  assign E6BEG0_input = {
    J2MID_GHb_END1,
    J2MID_EFb_END1,
    J2MID_CDb_END1,
    J2MID_ABb_END1,
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    SS4END0,
    E1END3,
    NN4END0
  };
  cus_mux161_buf inst_cus_mux161_buf_E6BEG0 (
      .A0 (E6BEG0_input[0]),
      .A1 (E6BEG0_input[1]),
      .A2 (E6BEG0_input[2]),
      .A3 (E6BEG0_input[3]),
      .A4 (E6BEG0_input[4]),
      .A5 (E6BEG0_input[5]),
      .A6 (E6BEG0_input[6]),
      .A7 (E6BEG0_input[7]),
      .A8 (E6BEG0_input[8]),
      .A9 (E6BEG0_input[9]),
      .A10(E6BEG0_input[10]),
      .A11(E6BEG0_input[11]),
      .A12(E6BEG0_input[12]),
      .A13(E6BEG0_input[13]),
      .A14(E6BEG0_input[14]),
      .A15(E6BEG0_input[15]),
      .S0 (ConfigBits[48+0]),
      .S0N(ConfigBits_N[48+0]),
      .S1 (ConfigBits[48+1]),
      .S1N(ConfigBits_N[48+1]),
      .S2 (ConfigBits[48+2]),
      .S2N(ConfigBits_N[48+2]),
      .S3 (ConfigBits[48+3]),
      .S3N(ConfigBits_N[48+3]),
      .X  (E6BEG0)
  );

  // switch matrix multiplexer  E6BEG1         MUX-16
  assign E6BEG1_input = {
    J2MID_GHa_END2,
    J2MID_EFa_END2,
    J2MID_CDa_END2,
    J2MID_ABa_END2,
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    SS4END3,
    E1END2,
    NN4END3
  };
  cus_mux161_buf inst_cus_mux161_buf_E6BEG1 (
      .A0 (E6BEG1_input[0]),
      .A1 (E6BEG1_input[1]),
      .A2 (E6BEG1_input[2]),
      .A3 (E6BEG1_input[3]),
      .A4 (E6BEG1_input[4]),
      .A5 (E6BEG1_input[5]),
      .A6 (E6BEG1_input[6]),
      .A7 (E6BEG1_input[7]),
      .A8 (E6BEG1_input[8]),
      .A9 (E6BEG1_input[9]),
      .A10(E6BEG1_input[10]),
      .A11(E6BEG1_input[11]),
      .A12(E6BEG1_input[12]),
      .A13(E6BEG1_input[13]),
      .A14(E6BEG1_input[14]),
      .A15(E6BEG1_input[15]),
      .S0 (ConfigBits[52+0]),
      .S0N(ConfigBits_N[52+0]),
      .S1 (ConfigBits[52+1]),
      .S1N(ConfigBits_N[52+1]),
      .S2 (ConfigBits[52+2]),
      .S2N(ConfigBits_N[52+2]),
      .S3 (ConfigBits[52+3]),
      .S3N(ConfigBits_N[52+3]),
      .X  (E6BEG1)
  );

  // switch matrix multiplexer  S1BEG0         MUX-4
  assign S1BEG0_input = {J_l_CD_END1, JE2END3, J2MID_CDb_END3, BD0};
  cus_mux41_buf inst_cus_mux41_buf_S1BEG0 (
      .A0 (S1BEG0_input[0]),
      .A1 (S1BEG0_input[1]),
      .A2 (S1BEG0_input[2]),
      .A3 (S1BEG0_input[3]),
      .S0 (ConfigBits[56+0]),
      .S0N(ConfigBits_N[56+0]),
      .S1 (ConfigBits[56+1]),
      .S1N(ConfigBits_N[56+1]),
      .X  (S1BEG0)
  );

  // switch matrix multiplexer  S1BEG1         MUX-4
  assign S1BEG1_input = {J_l_EF_END2, JE2END0, J2MID_EFb_END0, BD1};
  cus_mux41_buf inst_cus_mux41_buf_S1BEG1 (
      .A0 (S1BEG1_input[0]),
      .A1 (S1BEG1_input[1]),
      .A2 (S1BEG1_input[2]),
      .A3 (S1BEG1_input[3]),
      .S0 (ConfigBits[58+0]),
      .S0N(ConfigBits_N[58+0]),
      .S1 (ConfigBits[58+1]),
      .S1N(ConfigBits_N[58+1]),
      .X  (S1BEG1)
  );

  // switch matrix multiplexer  S1BEG2         MUX-4
  assign S1BEG2_input = {J_l_GH_END3, JE2END1, J2MID_GHb_END1, BD2};
  cus_mux41_buf inst_cus_mux41_buf_S1BEG2 (
      .A0 (S1BEG2_input[0]),
      .A1 (S1BEG2_input[1]),
      .A2 (S1BEG2_input[2]),
      .A3 (S1BEG2_input[3]),
      .S0 (ConfigBits[60+0]),
      .S0N(ConfigBits_N[60+0]),
      .S1 (ConfigBits[60+1]),
      .S1N(ConfigBits_N[60+1]),
      .X  (S1BEG2)
  );

  // switch matrix multiplexer  S1BEG3         MUX-4
  assign S1BEG3_input = {J_l_AB_END0, JE2END2, J2MID_ABb_END2, BD3};
  cus_mux41_buf inst_cus_mux41_buf_S1BEG3 (
      .A0 (S1BEG3_input[0]),
      .A1 (S1BEG3_input[1]),
      .A2 (S1BEG3_input[2]),
      .A3 (S1BEG3_input[3]),
      .S0 (ConfigBits[62+0]),
      .S0N(ConfigBits_N[62+0]),
      .S1 (ConfigBits[62+1]),
      .S1N(ConfigBits_N[62+1]),
      .X  (S1BEG3)
  );

  // switch matrix multiplexer  S2BEG0         MUX-1
  assign S2BEG0 = JS2END0;
  // switch matrix multiplexer  S2BEG1         MUX-1
  assign S2BEG1 = JS2END1;
  // switch matrix multiplexer  S2BEG2         MUX-1
  assign S2BEG2 = JS2END2;
  // switch matrix multiplexer  S2BEG3         MUX-1
  assign S2BEG3 = JS2END3;
  // switch matrix multiplexer  S2BEG4         MUX-1
  assign S2BEG4 = JS2END4;
  // switch matrix multiplexer  S2BEG5         MUX-1
  assign S2BEG5 = JS2END5;
  // switch matrix multiplexer  S2BEG6         MUX-1
  assign S2BEG6 = JS2END6;
  // switch matrix multiplexer  S2BEG7         MUX-1
  assign S2BEG7 = JS2END7;
  // switch matrix multiplexer  S2BEGb0         MUX-1
  assign S2BEGb0 = S2MID0;
  // switch matrix multiplexer  S2BEGb1         MUX-1
  assign S2BEGb1 = S2MID1;
  // switch matrix multiplexer  S2BEGb2         MUX-1
  assign S2BEGb2 = S2MID2;
  // switch matrix multiplexer  S2BEGb3         MUX-1
  assign S2BEGb3 = S2MID3;
  // switch matrix multiplexer  S2BEGb4         MUX-1
  assign S2BEGb4 = S2MID4;
  // switch matrix multiplexer  S2BEGb5         MUX-1
  assign S2BEGb5 = S2MID5;
  // switch matrix multiplexer  S2BEGb6         MUX-1
  assign S2BEGb6 = S2MID6;
  // switch matrix multiplexer  S2BEGb7         MUX-1
  assign S2BEGb7 = S2MID7;
  // switch matrix multiplexer  S4BEG0         MUX-4
  assign S4BEG0_input = {AD0, S4END1, S2END2, E6END1};
  cus_mux41_buf inst_cus_mux41_buf_S4BEG0 (
      .A0 (S4BEG0_input[0]),
      .A1 (S4BEG0_input[1]),
      .A2 (S4BEG0_input[2]),
      .A3 (S4BEG0_input[3]),
      .S0 (ConfigBits[64+0]),
      .S0N(ConfigBits_N[64+0]),
      .S1 (ConfigBits[64+1]),
      .S1N(ConfigBits_N[64+1]),
      .X  (S4BEG0)
  );

  // switch matrix multiplexer  S4BEG1         MUX-4
  assign S4BEG1_input = {AD1, S4END2, S2END3, E6END0};
  cus_mux41_buf inst_cus_mux41_buf_S4BEG1 (
      .A0 (S4BEG1_input[0]),
      .A1 (S4BEG1_input[1]),
      .A2 (S4BEG1_input[2]),
      .A3 (S4BEG1_input[3]),
      .S0 (ConfigBits[66+0]),
      .S0N(ConfigBits_N[66+0]),
      .S1 (ConfigBits[66+1]),
      .S1N(ConfigBits_N[66+1]),
      .X  (S4BEG1)
  );

  // switch matrix multiplexer  S4BEG2         MUX-4
  assign S4BEG2_input = {AD2, W6END1, S4END3, S2END0};
  cus_mux41_buf inst_cus_mux41_buf_S4BEG2 (
      .A0 (S4BEG2_input[0]),
      .A1 (S4BEG2_input[1]),
      .A2 (S4BEG2_input[2]),
      .A3 (S4BEG2_input[3]),
      .S0 (ConfigBits[68+0]),
      .S0N(ConfigBits_N[68+0]),
      .S1 (ConfigBits[68+1]),
      .S1N(ConfigBits_N[68+1]),
      .X  (S4BEG2)
  );

  // switch matrix multiplexer  S4BEG3         MUX-4
  assign S4BEG3_input = {AD3, W6END0, S4END0, S2END1};
  cus_mux41_buf inst_cus_mux41_buf_S4BEG3 (
      .A0 (S4BEG3_input[0]),
      .A1 (S4BEG3_input[1]),
      .A2 (S4BEG3_input[2]),
      .A3 (S4BEG3_input[3]),
      .S0 (ConfigBits[70+0]),
      .S0N(ConfigBits_N[70+0]),
      .S1 (ConfigBits[70+1]),
      .S1N(ConfigBits_N[70+1]),
      .X  (S4BEG3)
  );

  // switch matrix multiplexer  SS4BEG0         MUX-8
  assign SS4BEG0_input = {
    J2END_GH_END3, J2MID_CDb_END1, J2MID_ABb_END1, BD1, AD1, W1END2, E1END2, N1END2
  };
  cus_mux81_buf inst_cus_mux81_buf_SS4BEG0 (
      .A0 (SS4BEG0_input[0]),
      .A1 (SS4BEG0_input[1]),
      .A2 (SS4BEG0_input[2]),
      .A3 (SS4BEG0_input[3]),
      .A4 (SS4BEG0_input[4]),
      .A5 (SS4BEG0_input[5]),
      .A6 (SS4BEG0_input[6]),
      .A7 (SS4BEG0_input[7]),
      .S0 (ConfigBits[72+0]),
      .S0N(ConfigBits_N[72+0]),
      .S1 (ConfigBits[72+1]),
      .S1N(ConfigBits_N[72+1]),
      .S2 (ConfigBits[72+2]),
      .S2N(ConfigBits_N[72+2]),
      .X  (SS4BEG0)
  );

  // switch matrix multiplexer  SS4BEG1         MUX-8
  assign SS4BEG1_input = {
    J2END_EF_END3, J2MID_CDa_END2, J2MID_ABa_END2, BD2, AD2, W1END3, E1END3, N1END3
  };
  cus_mux81_buf inst_cus_mux81_buf_SS4BEG1 (
      .A0 (SS4BEG1_input[0]),
      .A1 (SS4BEG1_input[1]),
      .A2 (SS4BEG1_input[2]),
      .A3 (SS4BEG1_input[3]),
      .A4 (SS4BEG1_input[4]),
      .A5 (SS4BEG1_input[5]),
      .A6 (SS4BEG1_input[6]),
      .A7 (SS4BEG1_input[7]),
      .S0 (ConfigBits[75+0]),
      .S0N(ConfigBits_N[75+0]),
      .S1 (ConfigBits[75+1]),
      .S1N(ConfigBits_N[75+1]),
      .S2 (ConfigBits[75+2]),
      .S2N(ConfigBits_N[75+2]),
      .X  (SS4BEG1)
  );

  // switch matrix multiplexer  SS4BEG2         MUX-8
  assign SS4BEG2_input = {
    J2END_CD_END3, J2MID_GHb_END1, J2MID_EFb_END1, BD3, AD3, W1END0, E1END0, N1END0
  };
  cus_mux81_buf inst_cus_mux81_buf_SS4BEG2 (
      .A0 (SS4BEG2_input[0]),
      .A1 (SS4BEG2_input[1]),
      .A2 (SS4BEG2_input[2]),
      .A3 (SS4BEG2_input[3]),
      .A4 (SS4BEG2_input[4]),
      .A5 (SS4BEG2_input[5]),
      .A6 (SS4BEG2_input[6]),
      .A7 (SS4BEG2_input[7]),
      .S0 (ConfigBits[78+0]),
      .S0N(ConfigBits_N[78+0]),
      .S1 (ConfigBits[78+1]),
      .S1N(ConfigBits_N[78+1]),
      .S2 (ConfigBits[78+2]),
      .S2N(ConfigBits_N[78+2]),
      .X  (SS4BEG2)
  );

  // switch matrix multiplexer  SS4BEG3         MUX-8
  assign SS4BEG3_input = {
    J2END_AB_END3, J2MID_GHa_END2, J2MID_EFa_END2, BD0, AD0, W1END1, E1END1, N1END1
  };
  cus_mux81_buf inst_cus_mux81_buf_SS4BEG3 (
      .A0 (SS4BEG3_input[0]),
      .A1 (SS4BEG3_input[1]),
      .A2 (SS4BEG3_input[2]),
      .A3 (SS4BEG3_input[3]),
      .A4 (SS4BEG3_input[4]),
      .A5 (SS4BEG3_input[5]),
      .A6 (SS4BEG3_input[6]),
      .A7 (SS4BEG3_input[7]),
      .S0 (ConfigBits[81+0]),
      .S0N(ConfigBits_N[81+0]),
      .S1 (ConfigBits[81+1]),
      .S1N(ConfigBits_N[81+1]),
      .S2 (ConfigBits[81+2]),
      .S2N(ConfigBits_N[81+2]),
      .X  (SS4BEG3)
  );

  // switch matrix multiplexer  W1BEG0         MUX-4
  assign W1BEG0_input = {J_l_CD_END1, JS2END3, J2MID_CDb_END3, BD1};
  cus_mux41_buf inst_cus_mux41_buf_W1BEG0 (
      .A0 (W1BEG0_input[0]),
      .A1 (W1BEG0_input[1]),
      .A2 (W1BEG0_input[2]),
      .A3 (W1BEG0_input[3]),
      .S0 (ConfigBits[84+0]),
      .S0N(ConfigBits_N[84+0]),
      .S1 (ConfigBits[84+1]),
      .S1N(ConfigBits_N[84+1]),
      .X  (W1BEG0)
  );

  // switch matrix multiplexer  W1BEG1         MUX-4
  assign W1BEG1_input = {J_l_EF_END2, JS2END0, J2MID_EFb_END0, BD2};
  cus_mux41_buf inst_cus_mux41_buf_W1BEG1 (
      .A0 (W1BEG1_input[0]),
      .A1 (W1BEG1_input[1]),
      .A2 (W1BEG1_input[2]),
      .A3 (W1BEG1_input[3]),
      .S0 (ConfigBits[86+0]),
      .S0N(ConfigBits_N[86+0]),
      .S1 (ConfigBits[86+1]),
      .S1N(ConfigBits_N[86+1]),
      .X  (W1BEG1)
  );

  // switch matrix multiplexer  W1BEG2         MUX-4
  assign W1BEG2_input = {J_l_GH_END3, JS2END1, J2MID_GHb_END1, BD3};
  cus_mux41_buf inst_cus_mux41_buf_W1BEG2 (
      .A0 (W1BEG2_input[0]),
      .A1 (W1BEG2_input[1]),
      .A2 (W1BEG2_input[2]),
      .A3 (W1BEG2_input[3]),
      .S0 (ConfigBits[88+0]),
      .S0N(ConfigBits_N[88+0]),
      .S1 (ConfigBits[88+1]),
      .S1N(ConfigBits_N[88+1]),
      .X  (W1BEG2)
  );

  // switch matrix multiplexer  W1BEG3         MUX-4
  assign W1BEG3_input = {J_l_AB_END0, JS2END2, J2MID_ABb_END2, AD0};
  cus_mux41_buf inst_cus_mux41_buf_W1BEG3 (
      .A0 (W1BEG3_input[0]),
      .A1 (W1BEG3_input[1]),
      .A2 (W1BEG3_input[2]),
      .A3 (W1BEG3_input[3]),
      .S0 (ConfigBits[90+0]),
      .S0N(ConfigBits_N[90+0]),
      .S1 (ConfigBits[90+1]),
      .S1N(ConfigBits_N[90+1]),
      .X  (W1BEG3)
  );

  // switch matrix multiplexer  W2BEG0         MUX-1
  assign W2BEG0 = JW2END0;
  // switch matrix multiplexer  W2BEG1         MUX-1
  assign W2BEG1 = JW2END1;
  // switch matrix multiplexer  W2BEG2         MUX-1
  assign W2BEG2 = JW2END2;
  // switch matrix multiplexer  W2BEG3         MUX-1
  assign W2BEG3 = JW2END3;
  // switch matrix multiplexer  W2BEG4         MUX-1
  assign W2BEG4 = JW2END4;
  // switch matrix multiplexer  W2BEG5         MUX-1
  assign W2BEG5 = JW2END5;
  // switch matrix multiplexer  W2BEG6         MUX-1
  assign W2BEG6 = JW2END6;
  // switch matrix multiplexer  W2BEG7         MUX-1
  assign W2BEG7 = JW2END7;
  // switch matrix multiplexer  W2BEGb0         MUX-1
  assign W2BEGb0 = W2MID0;
  // switch matrix multiplexer  W2BEGb1         MUX-1
  assign W2BEGb1 = W2MID1;
  // switch matrix multiplexer  W2BEGb2         MUX-1
  assign W2BEGb2 = W2MID2;
  // switch matrix multiplexer  W2BEGb3         MUX-1
  assign W2BEGb3 = W2MID3;
  // switch matrix multiplexer  W2BEGb4         MUX-1
  assign W2BEGb4 = W2MID4;
  // switch matrix multiplexer  W2BEGb5         MUX-1
  assign W2BEGb5 = W2MID5;
  // switch matrix multiplexer  W2BEGb6         MUX-1
  assign W2BEGb6 = W2MID6;
  // switch matrix multiplexer  W2BEGb7         MUX-1
  assign W2BEGb7 = W2MID7;
  // switch matrix multiplexer  WW4BEG0         MUX-8
  assign WW4BEG0_input = {
    J2END_GH_END2, J2MID_CDb_END1, J2MID_ABb_END1, BD1, AD1, W1END2, S1END2, N1END2
  };
  cus_mux81_buf inst_cus_mux81_buf_WW4BEG0 (
      .A0 (WW4BEG0_input[0]),
      .A1 (WW4BEG0_input[1]),
      .A2 (WW4BEG0_input[2]),
      .A3 (WW4BEG0_input[3]),
      .A4 (WW4BEG0_input[4]),
      .A5 (WW4BEG0_input[5]),
      .A6 (WW4BEG0_input[6]),
      .A7 (WW4BEG0_input[7]),
      .S0 (ConfigBits[92+0]),
      .S0N(ConfigBits_N[92+0]),
      .S1 (ConfigBits[92+1]),
      .S1N(ConfigBits_N[92+1]),
      .S2 (ConfigBits[92+2]),
      .S2N(ConfigBits_N[92+2]),
      .X  (WW4BEG0)
  );

  // switch matrix multiplexer  WW4BEG1         MUX-8
  assign WW4BEG1_input = {
    J2END_EF_END2, J2MID_CDa_END2, J2MID_ABa_END2, BD2, AD2, W1END3, S1END3, N1END3
  };
  cus_mux81_buf inst_cus_mux81_buf_WW4BEG1 (
      .A0 (WW4BEG1_input[0]),
      .A1 (WW4BEG1_input[1]),
      .A2 (WW4BEG1_input[2]),
      .A3 (WW4BEG1_input[3]),
      .A4 (WW4BEG1_input[4]),
      .A5 (WW4BEG1_input[5]),
      .A6 (WW4BEG1_input[6]),
      .A7 (WW4BEG1_input[7]),
      .S0 (ConfigBits[95+0]),
      .S0N(ConfigBits_N[95+0]),
      .S1 (ConfigBits[95+1]),
      .S1N(ConfigBits_N[95+1]),
      .S2 (ConfigBits[95+2]),
      .S2N(ConfigBits_N[95+2]),
      .X  (WW4BEG1)
  );

  // switch matrix multiplexer  WW4BEG2         MUX-8
  assign WW4BEG2_input = {
    J2END_CD_END2, J2MID_GHb_END1, J2MID_EFb_END1, BD3, AD3, W1END0, S1END0, N1END0
  };
  cus_mux81_buf inst_cus_mux81_buf_WW4BEG2 (
      .A0 (WW4BEG2_input[0]),
      .A1 (WW4BEG2_input[1]),
      .A2 (WW4BEG2_input[2]),
      .A3 (WW4BEG2_input[3]),
      .A4 (WW4BEG2_input[4]),
      .A5 (WW4BEG2_input[5]),
      .A6 (WW4BEG2_input[6]),
      .A7 (WW4BEG2_input[7]),
      .S0 (ConfigBits[98+0]),
      .S0N(ConfigBits_N[98+0]),
      .S1 (ConfigBits[98+1]),
      .S1N(ConfigBits_N[98+1]),
      .S2 (ConfigBits[98+2]),
      .S2N(ConfigBits_N[98+2]),
      .X  (WW4BEG2)
  );

  // switch matrix multiplexer  WW4BEG3         MUX-8
  assign WW4BEG3_input = {
    J2END_AB_END2, J2MID_GHa_END2, J2MID_EFa_END2, BD0, AD0, W1END1, S1END1, N1END1
  };
  cus_mux81_buf inst_cus_mux81_buf_WW4BEG3 (
      .A0 (WW4BEG3_input[0]),
      .A1 (WW4BEG3_input[1]),
      .A2 (WW4BEG3_input[2]),
      .A3 (WW4BEG3_input[3]),
      .A4 (WW4BEG3_input[4]),
      .A5 (WW4BEG3_input[5]),
      .A6 (WW4BEG3_input[6]),
      .A7 (WW4BEG3_input[7]),
      .S0 (ConfigBits[101+0]),
      .S0N(ConfigBits_N[101+0]),
      .S1 (ConfigBits[101+1]),
      .S1N(ConfigBits_N[101+1]),
      .S2 (ConfigBits[101+2]),
      .S2N(ConfigBits_N[101+2]),
      .X  (WW4BEG3)
  );

  // switch matrix multiplexer  W6BEG0         MUX-16
  assign W6BEG0_input = {
    J2MID_GHb_END1,
    J2MID_EFb_END1,
    J2MID_CDb_END1,
    J2MID_ABb_END1,
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    SS4END1,
    E1END3,
    NN4END1
  };
  cus_mux161_buf inst_cus_mux161_buf_W6BEG0 (
      .A0 (W6BEG0_input[0]),
      .A1 (W6BEG0_input[1]),
      .A2 (W6BEG0_input[2]),
      .A3 (W6BEG0_input[3]),
      .A4 (W6BEG0_input[4]),
      .A5 (W6BEG0_input[5]),
      .A6 (W6BEG0_input[6]),
      .A7 (W6BEG0_input[7]),
      .A8 (W6BEG0_input[8]),
      .A9 (W6BEG0_input[9]),
      .A10(W6BEG0_input[10]),
      .A11(W6BEG0_input[11]),
      .A12(W6BEG0_input[12]),
      .A13(W6BEG0_input[13]),
      .A14(W6BEG0_input[14]),
      .A15(W6BEG0_input[15]),
      .S0 (ConfigBits[104+0]),
      .S0N(ConfigBits_N[104+0]),
      .S1 (ConfigBits[104+1]),
      .S1N(ConfigBits_N[104+1]),
      .S2 (ConfigBits[104+2]),
      .S2N(ConfigBits_N[104+2]),
      .S3 (ConfigBits[104+3]),
      .S3N(ConfigBits_N[104+3]),
      .X  (W6BEG0)
  );

  // switch matrix multiplexer  W6BEG1         MUX-16
  assign W6BEG1_input = {
    J2MID_GHa_END2,
    J2MID_EFa_END2,
    J2MID_CDa_END2,
    J2MID_ABa_END2,
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    SS4END2,
    E1END2,
    NN4END2
  };
  cus_mux161_buf inst_cus_mux161_buf_W6BEG1 (
      .A0 (W6BEG1_input[0]),
      .A1 (W6BEG1_input[1]),
      .A2 (W6BEG1_input[2]),
      .A3 (W6BEG1_input[3]),
      .A4 (W6BEG1_input[4]),
      .A5 (W6BEG1_input[5]),
      .A6 (W6BEG1_input[6]),
      .A7 (W6BEG1_input[7]),
      .A8 (W6BEG1_input[8]),
      .A9 (W6BEG1_input[9]),
      .A10(W6BEG1_input[10]),
      .A11(W6BEG1_input[11]),
      .A12(W6BEG1_input[12]),
      .A13(W6BEG1_input[13]),
      .A14(W6BEG1_input[14]),
      .A15(W6BEG1_input[15]),
      .S0 (ConfigBits[108+0]),
      .S0N(ConfigBits_N[108+0]),
      .S1 (ConfigBits[108+1]),
      .S1N(ConfigBits_N[108+1]),
      .S2 (ConfigBits[108+2]),
      .S2N(ConfigBits_N[108+2]),
      .S3 (ConfigBits[108+3]),
      .S3N(ConfigBits_N[108+3]),
      .X  (W6BEG1)
  );

  // switch matrix multiplexer  D0         MUX-4
  assign D0_input = {J_l_AB_END0, J2END_AB_END0, J2MID_ABb_END0, J2MID_ABa_END0};
  cus_mux41_buf inst_cus_mux41_buf_D0 (
      .A0 (D0_input[0]),
      .A1 (D0_input[1]),
      .A2 (D0_input[2]),
      .A3 (D0_input[3]),
      .S0 (ConfigBits[112+0]),
      .S0N(ConfigBits_N[112+0]),
      .S1 (ConfigBits[112+1]),
      .S1N(ConfigBits_N[112+1]),
      .X  (D0)
  );

  // switch matrix multiplexer  D1         MUX-4
  assign D1_input = {J_l_AB_END1, J2END_AB_END1, J2MID_ABb_END1, J2MID_ABa_END1};
  cus_mux41_buf inst_cus_mux41_buf_D1 (
      .A0 (D1_input[0]),
      .A1 (D1_input[1]),
      .A2 (D1_input[2]),
      .A3 (D1_input[3]),
      .S0 (ConfigBits[114+0]),
      .S0N(ConfigBits_N[114+0]),
      .S1 (ConfigBits[114+1]),
      .S1N(ConfigBits_N[114+1]),
      .X  (D1)
  );

  // switch matrix multiplexer  D2         MUX-4
  assign D2_input = {J_l_AB_END2, J2END_AB_END2, J2MID_ABb_END2, J2MID_ABa_END2};
  cus_mux41_buf inst_cus_mux41_buf_D2 (
      .A0 (D2_input[0]),
      .A1 (D2_input[1]),
      .A2 (D2_input[2]),
      .A3 (D2_input[3]),
      .S0 (ConfigBits[116+0]),
      .S0N(ConfigBits_N[116+0]),
      .S1 (ConfigBits[116+1]),
      .S1N(ConfigBits_N[116+1]),
      .X  (D2)
  );

  // switch matrix multiplexer  D3         MUX-4
  assign D3_input = {J_l_AB_END3, J2END_AB_END3, J2MID_ABb_END3, J2MID_ABa_END3};
  cus_mux41_buf inst_cus_mux41_buf_D3 (
      .A0 (D3_input[0]),
      .A1 (D3_input[1]),
      .A2 (D3_input[2]),
      .A3 (D3_input[3]),
      .S0 (ConfigBits[118+0]),
      .S0N(ConfigBits_N[118+0]),
      .S1 (ConfigBits[118+1]),
      .S1N(ConfigBits_N[118+1]),
      .X  (D3)
  );

  // switch matrix multiplexer  W_ADR0         MUX-4
  assign W_ADR0_input = {J_l_CD_END0, J2END_CD_END0, J2MID_CDb_END0, J2MID_CDa_END0};
  cus_mux41_buf inst_cus_mux41_buf_W_ADR0 (
      .A0 (W_ADR0_input[0]),
      .A1 (W_ADR0_input[1]),
      .A2 (W_ADR0_input[2]),
      .A3 (W_ADR0_input[3]),
      .S0 (ConfigBits[120+0]),
      .S0N(ConfigBits_N[120+0]),
      .S1 (ConfigBits[120+1]),
      .S1N(ConfigBits_N[120+1]),
      .X  (W_ADR0)
  );

  // switch matrix multiplexer  W_ADR1         MUX-4
  assign W_ADR1_input = {J_l_CD_END1, J2END_CD_END1, J2MID_CDb_END1, J2MID_CDa_END1};
  cus_mux41_buf inst_cus_mux41_buf_W_ADR1 (
      .A0 (W_ADR1_input[0]),
      .A1 (W_ADR1_input[1]),
      .A2 (W_ADR1_input[2]),
      .A3 (W_ADR1_input[3]),
      .S0 (ConfigBits[122+0]),
      .S0N(ConfigBits_N[122+0]),
      .S1 (ConfigBits[122+1]),
      .S1N(ConfigBits_N[122+1]),
      .X  (W_ADR1)
  );

  // switch matrix multiplexer  W_ADR2         MUX-4
  assign W_ADR2_input = {J_l_CD_END2, J2END_CD_END2, J2MID_CDb_END2, J2MID_CDa_END2};
  cus_mux41_buf inst_cus_mux41_buf_W_ADR2 (
      .A0 (W_ADR2_input[0]),
      .A1 (W_ADR2_input[1]),
      .A2 (W_ADR2_input[2]),
      .A3 (W_ADR2_input[3]),
      .S0 (ConfigBits[124+0]),
      .S0N(ConfigBits_N[124+0]),
      .S1 (ConfigBits[124+1]),
      .S1N(ConfigBits_N[124+1]),
      .X  (W_ADR2)
  );

  // switch matrix multiplexer  W_ADR3         MUX-4
  assign W_ADR3_input = {J_l_CD_END3, J2END_CD_END3, J2MID_CDb_END3, J2MID_CDa_END3};
  cus_mux41_buf inst_cus_mux41_buf_W_ADR3 (
      .A0 (W_ADR3_input[0]),
      .A1 (W_ADR3_input[1]),
      .A2 (W_ADR3_input[2]),
      .A3 (W_ADR3_input[3]),
      .S0 (ConfigBits[126+0]),
      .S0N(ConfigBits_N[126+0]),
      .S1 (ConfigBits[126+1]),
      .S1N(ConfigBits_N[126+1]),
      .X  (W_ADR3)
  );

  // switch matrix multiplexer  W_ADR4         MUX-8
  assign W_ADR4_input = {
    JW2END7, JS2END7, JN2END7, J2END_AB_END3, J2MID_EFb_END2, J2MID_EFa_END1, S2END0, N2END0
  };
  cus_mux81_buf inst_cus_mux81_buf_W_ADR4 (
      .A0 (W_ADR4_input[0]),
      .A1 (W_ADR4_input[1]),
      .A2 (W_ADR4_input[2]),
      .A3 (W_ADR4_input[3]),
      .A4 (W_ADR4_input[4]),
      .A5 (W_ADR4_input[5]),
      .A6 (W_ADR4_input[6]),
      .A7 (W_ADR4_input[7]),
      .S0 (ConfigBits[128+0]),
      .S0N(ConfigBits_N[128+0]),
      .S1 (ConfigBits[128+1]),
      .S1N(ConfigBits_N[128+1]),
      .S2 (ConfigBits[128+2]),
      .S2N(ConfigBits_N[128+2]),
      .X  (W_ADR4)
  );

  // switch matrix multiplexer  W_en         MUX-8
  assign W_en_input = {
    JW2END0, JS2END0, JN2END0, J2END_GH_END3, J2MID_CDb_END2, J2MID_CDa_END1, S2END3, N2END3
  };
  cus_mux81_buf inst_cus_mux81_buf_W_en (
      .A0 (W_en_input[0]),
      .A1 (W_en_input[1]),
      .A2 (W_en_input[2]),
      .A3 (W_en_input[3]),
      .A4 (W_en_input[4]),
      .A5 (W_en_input[5]),
      .A6 (W_en_input[6]),
      .A7 (W_en_input[7]),
      .S0 (ConfigBits[131+0]),
      .S0N(ConfigBits_N[131+0]),
      .S1 (ConfigBits[131+1]),
      .S1N(ConfigBits_N[131+1]),
      .S2 (ConfigBits[131+2]),
      .S2N(ConfigBits_N[131+2]),
      .X  (W_en)
  );

  // switch matrix multiplexer  A_ADR0         MUX-4
  assign A_ADR0_input = {J_l_EF_END0, J2END_EF_END0, J2MID_EFb_END0, J2MID_EFa_END0};
  cus_mux41_buf inst_cus_mux41_buf_A_ADR0 (
      .A0 (A_ADR0_input[0]),
      .A1 (A_ADR0_input[1]),
      .A2 (A_ADR0_input[2]),
      .A3 (A_ADR0_input[3]),
      .S0 (ConfigBits[134+0]),
      .S0N(ConfigBits_N[134+0]),
      .S1 (ConfigBits[134+1]),
      .S1N(ConfigBits_N[134+1]),
      .X  (A_ADR0)
  );

  // switch matrix multiplexer  A_ADR1         MUX-4
  assign A_ADR1_input = {J_l_EF_END1, J2END_EF_END1, J2MID_EFb_END1, J2MID_EFa_END1};
  cus_mux41_buf inst_cus_mux41_buf_A_ADR1 (
      .A0 (A_ADR1_input[0]),
      .A1 (A_ADR1_input[1]),
      .A2 (A_ADR1_input[2]),
      .A3 (A_ADR1_input[3]),
      .S0 (ConfigBits[136+0]),
      .S0N(ConfigBits_N[136+0]),
      .S1 (ConfigBits[136+1]),
      .S1N(ConfigBits_N[136+1]),
      .X  (A_ADR1)
  );

  // switch matrix multiplexer  A_ADR2         MUX-4
  assign A_ADR2_input = {J_l_EF_END2, J2END_EF_END2, J2MID_EFb_END2, J2MID_EFa_END2};
  cus_mux41_buf inst_cus_mux41_buf_A_ADR2 (
      .A0 (A_ADR2_input[0]),
      .A1 (A_ADR2_input[1]),
      .A2 (A_ADR2_input[2]),
      .A3 (A_ADR2_input[3]),
      .S0 (ConfigBits[138+0]),
      .S0N(ConfigBits_N[138+0]),
      .S1 (ConfigBits[138+1]),
      .S1N(ConfigBits_N[138+1]),
      .X  (A_ADR2)
  );

  // switch matrix multiplexer  A_ADR3         MUX-4
  assign A_ADR3_input = {J_l_EF_END3, J2END_EF_END3, J2MID_EFb_END3, J2MID_EFa_END3};
  cus_mux41_buf inst_cus_mux41_buf_A_ADR3 (
      .A0 (A_ADR3_input[0]),
      .A1 (A_ADR3_input[1]),
      .A2 (A_ADR3_input[2]),
      .A3 (A_ADR3_input[3]),
      .S0 (ConfigBits[140+0]),
      .S0N(ConfigBits_N[140+0]),
      .S1 (ConfigBits[140+1]),
      .S1N(ConfigBits_N[140+1]),
      .X  (A_ADR3)
  );

  // switch matrix multiplexer  A_ADR4         MUX-8
  assign A_ADR4_input = {
    JW2END5, JS2END5, JN2END5, J2END_CD_END3, J2MID_GHb_END2, J2MID_GHa_END1, S2END1, N2END1
  };
  cus_mux81_buf inst_cus_mux81_buf_A_ADR4 (
      .A0 (A_ADR4_input[0]),
      .A1 (A_ADR4_input[1]),
      .A2 (A_ADR4_input[2]),
      .A3 (A_ADR4_input[3]),
      .A4 (A_ADR4_input[4]),
      .A5 (A_ADR4_input[5]),
      .A6 (A_ADR4_input[6]),
      .A7 (A_ADR4_input[7]),
      .S0 (ConfigBits[142+0]),
      .S0N(ConfigBits_N[142+0]),
      .S1 (ConfigBits[142+1]),
      .S1N(ConfigBits_N[142+1]),
      .S2 (ConfigBits[142+2]),
      .S2N(ConfigBits_N[142+2]),
      .X  (A_ADR4)
  );

  // switch matrix multiplexer  B_ADR0         MUX-4
  assign B_ADR0_input = {J_l_GH_END0, J2END_GH_END0, J2MID_GHb_END0, J2MID_GHa_END0};
  cus_mux41_buf inst_cus_mux41_buf_B_ADR0 (
      .A0 (B_ADR0_input[0]),
      .A1 (B_ADR0_input[1]),
      .A2 (B_ADR0_input[2]),
      .A3 (B_ADR0_input[3]),
      .S0 (ConfigBits[145+0]),
      .S0N(ConfigBits_N[145+0]),
      .S1 (ConfigBits[145+1]),
      .S1N(ConfigBits_N[145+1]),
      .X  (B_ADR0)
  );

  // switch matrix multiplexer  B_ADR1         MUX-4
  assign B_ADR1_input = {J_l_GH_END1, J2END_GH_END1, J2MID_GHb_END1, J2MID_GHa_END1};
  cus_mux41_buf inst_cus_mux41_buf_B_ADR1 (
      .A0 (B_ADR1_input[0]),
      .A1 (B_ADR1_input[1]),
      .A2 (B_ADR1_input[2]),
      .A3 (B_ADR1_input[3]),
      .S0 (ConfigBits[147+0]),
      .S0N(ConfigBits_N[147+0]),
      .S1 (ConfigBits[147+1]),
      .S1N(ConfigBits_N[147+1]),
      .X  (B_ADR1)
  );

  // switch matrix multiplexer  B_ADR2         MUX-4
  assign B_ADR2_input = {J_l_GH_END2, J2END_GH_END2, J2MID_GHb_END2, J2MID_GHa_END2};
  cus_mux41_buf inst_cus_mux41_buf_B_ADR2 (
      .A0 (B_ADR2_input[0]),
      .A1 (B_ADR2_input[1]),
      .A2 (B_ADR2_input[2]),
      .A3 (B_ADR2_input[3]),
      .S0 (ConfigBits[149+0]),
      .S0N(ConfigBits_N[149+0]),
      .S1 (ConfigBits[149+1]),
      .S1N(ConfigBits_N[149+1]),
      .X  (B_ADR2)
  );

  // switch matrix multiplexer  B_ADR3         MUX-4
  assign B_ADR3_input = {J_l_GH_END3, J2END_GH_END3, J2MID_GHb_END3, J2MID_GHa_END3};
  cus_mux41_buf inst_cus_mux41_buf_B_ADR3 (
      .A0 (B_ADR3_input[0]),
      .A1 (B_ADR3_input[1]),
      .A2 (B_ADR3_input[2]),
      .A3 (B_ADR3_input[3]),
      .S0 (ConfigBits[151+0]),
      .S0N(ConfigBits_N[151+0]),
      .S1 (ConfigBits[151+1]),
      .S1N(ConfigBits_N[151+1]),
      .X  (B_ADR3)
  );

  // switch matrix multiplexer  B_ADR4         MUX-8
  assign B_ADR4_input = {
    JW2END6, JS2END6, JN2END6, J2END_EF_END3, J2MID_ABb_END2, J2MID_ABa_END1, S2END2, N2END2
  };
  cus_mux81_buf inst_cus_mux81_buf_B_ADR4 (
      .A0 (B_ADR4_input[0]),
      .A1 (B_ADR4_input[1]),
      .A2 (B_ADR4_input[2]),
      .A3 (B_ADR4_input[3]),
      .A4 (B_ADR4_input[4]),
      .A5 (B_ADR4_input[5]),
      .A6 (B_ADR4_input[6]),
      .A7 (B_ADR4_input[7]),
      .S0 (ConfigBits[153+0]),
      .S0N(ConfigBits_N[153+0]),
      .S1 (ConfigBits[153+1]),
      .S1N(ConfigBits_N[153+1]),
      .S2 (ConfigBits[153+2]),
      .S2N(ConfigBits_N[153+2]),
      .X  (B_ADR4)
  );

  // switch matrix multiplexer  J2MID_ABa_BEG0         MUX-4
  assign J2MID_ABa_BEG0_input = {JN2END3, W2MID6, S2MID6, N2MID6};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG0 (
      .A0 (J2MID_ABa_BEG0_input[0]),
      .A1 (J2MID_ABa_BEG0_input[1]),
      .A2 (J2MID_ABa_BEG0_input[2]),
      .A3 (J2MID_ABa_BEG0_input[3]),
      .S0 (ConfigBits[156+0]),
      .S0N(ConfigBits_N[156+0]),
      .S1 (ConfigBits[156+1]),
      .S1N(ConfigBits_N[156+1]),
      .X  (J2MID_ABa_BEG0)
  );

  // switch matrix multiplexer  J2MID_ABa_BEG1         MUX-4
  assign J2MID_ABa_BEG1_input = {JE2END3, W2MID2, S2MID2, E2MID2};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG1 (
      .A0 (J2MID_ABa_BEG1_input[0]),
      .A1 (J2MID_ABa_BEG1_input[1]),
      .A2 (J2MID_ABa_BEG1_input[2]),
      .A3 (J2MID_ABa_BEG1_input[3]),
      .S0 (ConfigBits[158+0]),
      .S0N(ConfigBits_N[158+0]),
      .S1 (ConfigBits[158+1]),
      .S1N(ConfigBits_N[158+1]),
      .X  (J2MID_ABa_BEG1)
  );

  // switch matrix multiplexer  J2MID_ABa_BEG2         MUX-4
  assign J2MID_ABa_BEG2_input = {JS2END3, W2MID4, E2MID4, N2MID4};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG2 (
      .A0 (J2MID_ABa_BEG2_input[0]),
      .A1 (J2MID_ABa_BEG2_input[1]),
      .A2 (J2MID_ABa_BEG2_input[2]),
      .A3 (J2MID_ABa_BEG2_input[3]),
      .S0 (ConfigBits[160+0]),
      .S0N(ConfigBits_N[160+0]),
      .S1 (ConfigBits[160+1]),
      .S1N(ConfigBits_N[160+1]),
      .X  (J2MID_ABa_BEG2)
  );

  // switch matrix multiplexer  J2MID_ABa_BEG3         MUX-4
  assign J2MID_ABa_BEG3_input = {JW2END3, S2MID0, E2MID0, N2MID0};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG3 (
      .A0 (J2MID_ABa_BEG3_input[0]),
      .A1 (J2MID_ABa_BEG3_input[1]),
      .A2 (J2MID_ABa_BEG3_input[2]),
      .A3 (J2MID_ABa_BEG3_input[3]),
      .S0 (ConfigBits[162+0]),
      .S0N(ConfigBits_N[162+0]),
      .S1 (ConfigBits[162+1]),
      .S1N(ConfigBits_N[162+1]),
      .X  (J2MID_ABa_BEG3)
  );

  // switch matrix multiplexer  J2MID_CDa_BEG0         MUX-4
  assign J2MID_CDa_BEG0_input = {JN2END4, W2MID6, S2MID6, E2MID6};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG0 (
      .A0 (J2MID_CDa_BEG0_input[0]),
      .A1 (J2MID_CDa_BEG0_input[1]),
      .A2 (J2MID_CDa_BEG0_input[2]),
      .A3 (J2MID_CDa_BEG0_input[3]),
      .S0 (ConfigBits[164+0]),
      .S0N(ConfigBits_N[164+0]),
      .S1 (ConfigBits[164+1]),
      .S1N(ConfigBits_N[164+1]),
      .X  (J2MID_CDa_BEG0)
  );

  // switch matrix multiplexer  J2MID_CDa_BEG1         MUX-4
  assign J2MID_CDa_BEG1_input = {JE2END4, W2MID2, E2MID2, N2MID2};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG1 (
      .A0 (J2MID_CDa_BEG1_input[0]),
      .A1 (J2MID_CDa_BEG1_input[1]),
      .A2 (J2MID_CDa_BEG1_input[2]),
      .A3 (J2MID_CDa_BEG1_input[3]),
      .S0 (ConfigBits[166+0]),
      .S0N(ConfigBits_N[166+0]),
      .S1 (ConfigBits[166+1]),
      .S1N(ConfigBits_N[166+1]),
      .X  (J2MID_CDa_BEG1)
  );

  // switch matrix multiplexer  J2MID_CDa_BEG2         MUX-4
  assign J2MID_CDa_BEG2_input = {JS2END4, S2MID4, E2MID4, N2MID4};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG2 (
      .A0 (J2MID_CDa_BEG2_input[0]),
      .A1 (J2MID_CDa_BEG2_input[1]),
      .A2 (J2MID_CDa_BEG2_input[2]),
      .A3 (J2MID_CDa_BEG2_input[3]),
      .S0 (ConfigBits[168+0]),
      .S0N(ConfigBits_N[168+0]),
      .S1 (ConfigBits[168+1]),
      .S1N(ConfigBits_N[168+1]),
      .X  (J2MID_CDa_BEG2)
  );

  // switch matrix multiplexer  J2MID_CDa_BEG3         MUX-4
  assign J2MID_CDa_BEG3_input = {JW2END4, W2MID0, S2MID0, N2MID0};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG3 (
      .A0 (J2MID_CDa_BEG3_input[0]),
      .A1 (J2MID_CDa_BEG3_input[1]),
      .A2 (J2MID_CDa_BEG3_input[2]),
      .A3 (J2MID_CDa_BEG3_input[3]),
      .S0 (ConfigBits[170+0]),
      .S0N(ConfigBits_N[170+0]),
      .S1 (ConfigBits[170+1]),
      .S1N(ConfigBits_N[170+1]),
      .X  (J2MID_CDa_BEG3)
  );

  // switch matrix multiplexer  J2MID_EFa_BEG0         MUX-4
  assign J2MID_EFa_BEG0_input = {JN2END5, W2MID6, E2MID6, N2MID6};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG0 (
      .A0 (J2MID_EFa_BEG0_input[0]),
      .A1 (J2MID_EFa_BEG0_input[1]),
      .A2 (J2MID_EFa_BEG0_input[2]),
      .A3 (J2MID_EFa_BEG0_input[3]),
      .S0 (ConfigBits[172+0]),
      .S0N(ConfigBits_N[172+0]),
      .S1 (ConfigBits[172+1]),
      .S1N(ConfigBits_N[172+1]),
      .X  (J2MID_EFa_BEG0)
  );

  // switch matrix multiplexer  J2MID_EFa_BEG1         MUX-4
  assign J2MID_EFa_BEG1_input = {JE2END5, S2MID2, E2MID2, N2MID2};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG1 (
      .A0 (J2MID_EFa_BEG1_input[0]),
      .A1 (J2MID_EFa_BEG1_input[1]),
      .A2 (J2MID_EFa_BEG1_input[2]),
      .A3 (J2MID_EFa_BEG1_input[3]),
      .S0 (ConfigBits[174+0]),
      .S0N(ConfigBits_N[174+0]),
      .S1 (ConfigBits[174+1]),
      .S1N(ConfigBits_N[174+1]),
      .X  (J2MID_EFa_BEG1)
  );

  // switch matrix multiplexer  J2MID_EFa_BEG2         MUX-4
  assign J2MID_EFa_BEG2_input = {JS2END5, W2MID4, S2MID4, N2MID4};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG2 (
      .A0 (J2MID_EFa_BEG2_input[0]),
      .A1 (J2MID_EFa_BEG2_input[1]),
      .A2 (J2MID_EFa_BEG2_input[2]),
      .A3 (J2MID_EFa_BEG2_input[3]),
      .S0 (ConfigBits[176+0]),
      .S0N(ConfigBits_N[176+0]),
      .S1 (ConfigBits[176+1]),
      .S1N(ConfigBits_N[176+1]),
      .X  (J2MID_EFa_BEG2)
  );

  // switch matrix multiplexer  J2MID_EFa_BEG3         MUX-4
  assign J2MID_EFa_BEG3_input = {JW2END5, W2MID0, S2MID0, E2MID0};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG3 (
      .A0 (J2MID_EFa_BEG3_input[0]),
      .A1 (J2MID_EFa_BEG3_input[1]),
      .A2 (J2MID_EFa_BEG3_input[2]),
      .A3 (J2MID_EFa_BEG3_input[3]),
      .S0 (ConfigBits[178+0]),
      .S0N(ConfigBits_N[178+0]),
      .S1 (ConfigBits[178+1]),
      .S1N(ConfigBits_N[178+1]),
      .X  (J2MID_EFa_BEG3)
  );

  // switch matrix multiplexer  J2MID_GHa_BEG0         MUX-4
  assign J2MID_GHa_BEG0_input = {JN2END6, S2MID6, E2MID6, N2MID6};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG0 (
      .A0 (J2MID_GHa_BEG0_input[0]),
      .A1 (J2MID_GHa_BEG0_input[1]),
      .A2 (J2MID_GHa_BEG0_input[2]),
      .A3 (J2MID_GHa_BEG0_input[3]),
      .S0 (ConfigBits[180+0]),
      .S0N(ConfigBits_N[180+0]),
      .S1 (ConfigBits[180+1]),
      .S1N(ConfigBits_N[180+1]),
      .X  (J2MID_GHa_BEG0)
  );

  // switch matrix multiplexer  J2MID_GHa_BEG1         MUX-4
  assign J2MID_GHa_BEG1_input = {JE2END6, W2MID2, S2MID2, N2MID2};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG1 (
      .A0 (J2MID_GHa_BEG1_input[0]),
      .A1 (J2MID_GHa_BEG1_input[1]),
      .A2 (J2MID_GHa_BEG1_input[2]),
      .A3 (J2MID_GHa_BEG1_input[3]),
      .S0 (ConfigBits[182+0]),
      .S0N(ConfigBits_N[182+0]),
      .S1 (ConfigBits[182+1]),
      .S1N(ConfigBits_N[182+1]),
      .X  (J2MID_GHa_BEG1)
  );

  // switch matrix multiplexer  J2MID_GHa_BEG2         MUX-4
  assign J2MID_GHa_BEG2_input = {JS2END6, W2MID4, S2MID4, E2MID4};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG2 (
      .A0 (J2MID_GHa_BEG2_input[0]),
      .A1 (J2MID_GHa_BEG2_input[1]),
      .A2 (J2MID_GHa_BEG2_input[2]),
      .A3 (J2MID_GHa_BEG2_input[3]),
      .S0 (ConfigBits[184+0]),
      .S0N(ConfigBits_N[184+0]),
      .S1 (ConfigBits[184+1]),
      .S1N(ConfigBits_N[184+1]),
      .X  (J2MID_GHa_BEG2)
  );

  // switch matrix multiplexer  J2MID_GHa_BEG3         MUX-4
  assign J2MID_GHa_BEG3_input = {JW2END6, W2MID0, E2MID0, N2MID0};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG3 (
      .A0 (J2MID_GHa_BEG3_input[0]),
      .A1 (J2MID_GHa_BEG3_input[1]),
      .A2 (J2MID_GHa_BEG3_input[2]),
      .A3 (J2MID_GHa_BEG3_input[3]),
      .S0 (ConfigBits[186+0]),
      .S0N(ConfigBits_N[186+0]),
      .S1 (ConfigBits[186+1]),
      .S1N(ConfigBits_N[186+1]),
      .X  (J2MID_GHa_BEG3)
  );

  // switch matrix multiplexer  J2MID_ABb_BEG0         MUX-4
  assign J2MID_ABb_BEG0_input = {W2MID7, S2MID7, E2MID7, N2MID7};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG0 (
      .A0 (J2MID_ABb_BEG0_input[0]),
      .A1 (J2MID_ABb_BEG0_input[1]),
      .A2 (J2MID_ABb_BEG0_input[2]),
      .A3 (J2MID_ABb_BEG0_input[3]),
      .S0 (ConfigBits[188+0]),
      .S0N(ConfigBits_N[188+0]),
      .S1 (ConfigBits[188+1]),
      .S1N(ConfigBits_N[188+1]),
      .X  (J2MID_ABb_BEG0)
  );

  // switch matrix multiplexer  J2MID_ABb_BEG1         MUX-4
  assign J2MID_ABb_BEG1_input = {W2MID3, S2MID3, E2MID3, N2MID3};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG1 (
      .A0 (J2MID_ABb_BEG1_input[0]),
      .A1 (J2MID_ABb_BEG1_input[1]),
      .A2 (J2MID_ABb_BEG1_input[2]),
      .A3 (J2MID_ABb_BEG1_input[3]),
      .S0 (ConfigBits[190+0]),
      .S0N(ConfigBits_N[190+0]),
      .S1 (ConfigBits[190+1]),
      .S1N(ConfigBits_N[190+1]),
      .X  (J2MID_ABb_BEG1)
  );

  // switch matrix multiplexer  J2MID_ABb_BEG2         MUX-4
  assign J2MID_ABb_BEG2_input = {W2MID5, S2MID5, E2MID5, N2MID5};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG2 (
      .A0 (J2MID_ABb_BEG2_input[0]),
      .A1 (J2MID_ABb_BEG2_input[1]),
      .A2 (J2MID_ABb_BEG2_input[2]),
      .A3 (J2MID_ABb_BEG2_input[3]),
      .S0 (ConfigBits[192+0]),
      .S0N(ConfigBits_N[192+0]),
      .S1 (ConfigBits[192+1]),
      .S1N(ConfigBits_N[192+1]),
      .X  (J2MID_ABb_BEG2)
  );

  // switch matrix multiplexer  J2MID_ABb_BEG3         MUX-4
  assign J2MID_ABb_BEG3_input = {W2MID1, S2MID1, E2MID1, N2MID1};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG3 (
      .A0 (J2MID_ABb_BEG3_input[0]),
      .A1 (J2MID_ABb_BEG3_input[1]),
      .A2 (J2MID_ABb_BEG3_input[2]),
      .A3 (J2MID_ABb_BEG3_input[3]),
      .S0 (ConfigBits[194+0]),
      .S0N(ConfigBits_N[194+0]),
      .S1 (ConfigBits[194+1]),
      .S1N(ConfigBits_N[194+1]),
      .X  (J2MID_ABb_BEG3)
  );

  // switch matrix multiplexer  J2MID_CDb_BEG0         MUX-4
  assign J2MID_CDb_BEG0_input = {W2MID7, S2MID7, E2MID7, N2MID7};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG0 (
      .A0 (J2MID_CDb_BEG0_input[0]),
      .A1 (J2MID_CDb_BEG0_input[1]),
      .A2 (J2MID_CDb_BEG0_input[2]),
      .A3 (J2MID_CDb_BEG0_input[3]),
      .S0 (ConfigBits[196+0]),
      .S0N(ConfigBits_N[196+0]),
      .S1 (ConfigBits[196+1]),
      .S1N(ConfigBits_N[196+1]),
      .X  (J2MID_CDb_BEG0)
  );

  // switch matrix multiplexer  J2MID_CDb_BEG1         MUX-4
  assign J2MID_CDb_BEG1_input = {W2MID3, S2MID3, E2MID3, N2MID3};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG1 (
      .A0 (J2MID_CDb_BEG1_input[0]),
      .A1 (J2MID_CDb_BEG1_input[1]),
      .A2 (J2MID_CDb_BEG1_input[2]),
      .A3 (J2MID_CDb_BEG1_input[3]),
      .S0 (ConfigBits[198+0]),
      .S0N(ConfigBits_N[198+0]),
      .S1 (ConfigBits[198+1]),
      .S1N(ConfigBits_N[198+1]),
      .X  (J2MID_CDb_BEG1)
  );

  // switch matrix multiplexer  J2MID_CDb_BEG2         MUX-4
  assign J2MID_CDb_BEG2_input = {W2MID5, S2MID5, E2MID5, N2MID5};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG2 (
      .A0 (J2MID_CDb_BEG2_input[0]),
      .A1 (J2MID_CDb_BEG2_input[1]),
      .A2 (J2MID_CDb_BEG2_input[2]),
      .A3 (J2MID_CDb_BEG2_input[3]),
      .S0 (ConfigBits[200+0]),
      .S0N(ConfigBits_N[200+0]),
      .S1 (ConfigBits[200+1]),
      .S1N(ConfigBits_N[200+1]),
      .X  (J2MID_CDb_BEG2)
  );

  // switch matrix multiplexer  J2MID_CDb_BEG3         MUX-4
  assign J2MID_CDb_BEG3_input = {W2MID1, S2MID1, E2MID1, N2MID1};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG3 (
      .A0 (J2MID_CDb_BEG3_input[0]),
      .A1 (J2MID_CDb_BEG3_input[1]),
      .A2 (J2MID_CDb_BEG3_input[2]),
      .A3 (J2MID_CDb_BEG3_input[3]),
      .S0 (ConfigBits[202+0]),
      .S0N(ConfigBits_N[202+0]),
      .S1 (ConfigBits[202+1]),
      .S1N(ConfigBits_N[202+1]),
      .X  (J2MID_CDb_BEG3)
  );

  // switch matrix multiplexer  J2MID_EFb_BEG0         MUX-4
  assign J2MID_EFb_BEG0_input = {W2MID7, S2MID7, E2MID7, N2MID7};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG0 (
      .A0 (J2MID_EFb_BEG0_input[0]),
      .A1 (J2MID_EFb_BEG0_input[1]),
      .A2 (J2MID_EFb_BEG0_input[2]),
      .A3 (J2MID_EFb_BEG0_input[3]),
      .S0 (ConfigBits[204+0]),
      .S0N(ConfigBits_N[204+0]),
      .S1 (ConfigBits[204+1]),
      .S1N(ConfigBits_N[204+1]),
      .X  (J2MID_EFb_BEG0)
  );

  // switch matrix multiplexer  J2MID_EFb_BEG1         MUX-4
  assign J2MID_EFb_BEG1_input = {W2MID3, S2MID3, E2MID3, N2MID3};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG1 (
      .A0 (J2MID_EFb_BEG1_input[0]),
      .A1 (J2MID_EFb_BEG1_input[1]),
      .A2 (J2MID_EFb_BEG1_input[2]),
      .A3 (J2MID_EFb_BEG1_input[3]),
      .S0 (ConfigBits[206+0]),
      .S0N(ConfigBits_N[206+0]),
      .S1 (ConfigBits[206+1]),
      .S1N(ConfigBits_N[206+1]),
      .X  (J2MID_EFb_BEG1)
  );

  // switch matrix multiplexer  J2MID_EFb_BEG2         MUX-4
  assign J2MID_EFb_BEG2_input = {W2MID5, S2MID5, E2MID5, N2MID5};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG2 (
      .A0 (J2MID_EFb_BEG2_input[0]),
      .A1 (J2MID_EFb_BEG2_input[1]),
      .A2 (J2MID_EFb_BEG2_input[2]),
      .A3 (J2MID_EFb_BEG2_input[3]),
      .S0 (ConfigBits[208+0]),
      .S0N(ConfigBits_N[208+0]),
      .S1 (ConfigBits[208+1]),
      .S1N(ConfigBits_N[208+1]),
      .X  (J2MID_EFb_BEG2)
  );

  // switch matrix multiplexer  J2MID_EFb_BEG3         MUX-4
  assign J2MID_EFb_BEG3_input = {W2MID1, S2MID1, E2MID1, N2MID1};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG3 (
      .A0 (J2MID_EFb_BEG3_input[0]),
      .A1 (J2MID_EFb_BEG3_input[1]),
      .A2 (J2MID_EFb_BEG3_input[2]),
      .A3 (J2MID_EFb_BEG3_input[3]),
      .S0 (ConfigBits[210+0]),
      .S0N(ConfigBits_N[210+0]),
      .S1 (ConfigBits[210+1]),
      .S1N(ConfigBits_N[210+1]),
      .X  (J2MID_EFb_BEG3)
  );

  // switch matrix multiplexer  J2MID_GHb_BEG0         MUX-4
  assign J2MID_GHb_BEG0_input = {W2MID7, S2MID7, E2MID7, N2MID7};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG0 (
      .A0 (J2MID_GHb_BEG0_input[0]),
      .A1 (J2MID_GHb_BEG0_input[1]),
      .A2 (J2MID_GHb_BEG0_input[2]),
      .A3 (J2MID_GHb_BEG0_input[3]),
      .S0 (ConfigBits[212+0]),
      .S0N(ConfigBits_N[212+0]),
      .S1 (ConfigBits[212+1]),
      .S1N(ConfigBits_N[212+1]),
      .X  (J2MID_GHb_BEG0)
  );

  // switch matrix multiplexer  J2MID_GHb_BEG1         MUX-4
  assign J2MID_GHb_BEG1_input = {W2MID3, S2MID3, E2MID3, N2MID3};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG1 (
      .A0 (J2MID_GHb_BEG1_input[0]),
      .A1 (J2MID_GHb_BEG1_input[1]),
      .A2 (J2MID_GHb_BEG1_input[2]),
      .A3 (J2MID_GHb_BEG1_input[3]),
      .S0 (ConfigBits[214+0]),
      .S0N(ConfigBits_N[214+0]),
      .S1 (ConfigBits[214+1]),
      .S1N(ConfigBits_N[214+1]),
      .X  (J2MID_GHb_BEG1)
  );

  // switch matrix multiplexer  J2MID_GHb_BEG2         MUX-4
  assign J2MID_GHb_BEG2_input = {W2MID5, S2MID5, E2MID5, N2MID5};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG2 (
      .A0 (J2MID_GHb_BEG2_input[0]),
      .A1 (J2MID_GHb_BEG2_input[1]),
      .A2 (J2MID_GHb_BEG2_input[2]),
      .A3 (J2MID_GHb_BEG2_input[3]),
      .S0 (ConfigBits[216+0]),
      .S0N(ConfigBits_N[216+0]),
      .S1 (ConfigBits[216+1]),
      .S1N(ConfigBits_N[216+1]),
      .X  (J2MID_GHb_BEG2)
  );

  // switch matrix multiplexer  J2MID_GHb_BEG3         MUX-4
  assign J2MID_GHb_BEG3_input = {W2MID1, S2MID1, E2MID1, N2MID1};
  cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG3 (
      .A0 (J2MID_GHb_BEG3_input[0]),
      .A1 (J2MID_GHb_BEG3_input[1]),
      .A2 (J2MID_GHb_BEG3_input[2]),
      .A3 (J2MID_GHb_BEG3_input[3]),
      .S0 (ConfigBits[218+0]),
      .S0N(ConfigBits_N[218+0]),
      .S1 (ConfigBits[218+1]),
      .S1N(ConfigBits_N[218+1]),
      .X  (J2MID_GHb_BEG3)
  );

  // switch matrix multiplexer  J2END_AB_BEG0         MUX-4
  assign J2END_AB_BEG0_input = {W2END6, S2END6, E2END6, N2END6};
  cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG0 (
      .A0 (J2END_AB_BEG0_input[0]),
      .A1 (J2END_AB_BEG0_input[1]),
      .A2 (J2END_AB_BEG0_input[2]),
      .A3 (J2END_AB_BEG0_input[3]),
      .S0 (ConfigBits[220+0]),
      .S0N(ConfigBits_N[220+0]),
      .S1 (ConfigBits[220+1]),
      .S1N(ConfigBits_N[220+1]),
      .X  (J2END_AB_BEG0)
  );

  // switch matrix multiplexer  J2END_AB_BEG1         MUX-4
  assign J2END_AB_BEG1_input = {W2END2, S2END2, E2END2, N2END2};
  cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG1 (
      .A0 (J2END_AB_BEG1_input[0]),
      .A1 (J2END_AB_BEG1_input[1]),
      .A2 (J2END_AB_BEG1_input[2]),
      .A3 (J2END_AB_BEG1_input[3]),
      .S0 (ConfigBits[222+0]),
      .S0N(ConfigBits_N[222+0]),
      .S1 (ConfigBits[222+1]),
      .S1N(ConfigBits_N[222+1]),
      .X  (J2END_AB_BEG1)
  );

  // switch matrix multiplexer  J2END_AB_BEG2         MUX-4
  assign J2END_AB_BEG2_input = {W2END4, S2END4, E2END4, N2END4};
  cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG2 (
      .A0 (J2END_AB_BEG2_input[0]),
      .A1 (J2END_AB_BEG2_input[1]),
      .A2 (J2END_AB_BEG2_input[2]),
      .A3 (J2END_AB_BEG2_input[3]),
      .S0 (ConfigBits[224+0]),
      .S0N(ConfigBits_N[224+0]),
      .S1 (ConfigBits[224+1]),
      .S1N(ConfigBits_N[224+1]),
      .X  (J2END_AB_BEG2)
  );

  // switch matrix multiplexer  J2END_AB_BEG3         MUX-4
  assign J2END_AB_BEG3_input = {W2END0, S2END0, E2END0, N2END0};
  cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG3 (
      .A0 (J2END_AB_BEG3_input[0]),
      .A1 (J2END_AB_BEG3_input[1]),
      .A2 (J2END_AB_BEG3_input[2]),
      .A3 (J2END_AB_BEG3_input[3]),
      .S0 (ConfigBits[226+0]),
      .S0N(ConfigBits_N[226+0]),
      .S1 (ConfigBits[226+1]),
      .S1N(ConfigBits_N[226+1]),
      .X  (J2END_AB_BEG3)
  );

  // switch matrix multiplexer  J2END_CD_BEG0         MUX-4
  assign J2END_CD_BEG0_input = {W2END6, S2END6, E2END6, N2END6};
  cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG0 (
      .A0 (J2END_CD_BEG0_input[0]),
      .A1 (J2END_CD_BEG0_input[1]),
      .A2 (J2END_CD_BEG0_input[2]),
      .A3 (J2END_CD_BEG0_input[3]),
      .S0 (ConfigBits[228+0]),
      .S0N(ConfigBits_N[228+0]),
      .S1 (ConfigBits[228+1]),
      .S1N(ConfigBits_N[228+1]),
      .X  (J2END_CD_BEG0)
  );

  // switch matrix multiplexer  J2END_CD_BEG1         MUX-4
  assign J2END_CD_BEG1_input = {W2END2, S2END2, E2END2, N2END2};
  cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG1 (
      .A0 (J2END_CD_BEG1_input[0]),
      .A1 (J2END_CD_BEG1_input[1]),
      .A2 (J2END_CD_BEG1_input[2]),
      .A3 (J2END_CD_BEG1_input[3]),
      .S0 (ConfigBits[230+0]),
      .S0N(ConfigBits_N[230+0]),
      .S1 (ConfigBits[230+1]),
      .S1N(ConfigBits_N[230+1]),
      .X  (J2END_CD_BEG1)
  );

  // switch matrix multiplexer  J2END_CD_BEG2         MUX-4
  assign J2END_CD_BEG2_input = {W2END4, S2END4, E2END4, N2END4};
  cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG2 (
      .A0 (J2END_CD_BEG2_input[0]),
      .A1 (J2END_CD_BEG2_input[1]),
      .A2 (J2END_CD_BEG2_input[2]),
      .A3 (J2END_CD_BEG2_input[3]),
      .S0 (ConfigBits[232+0]),
      .S0N(ConfigBits_N[232+0]),
      .S1 (ConfigBits[232+1]),
      .S1N(ConfigBits_N[232+1]),
      .X  (J2END_CD_BEG2)
  );

  // switch matrix multiplexer  J2END_CD_BEG3         MUX-4
  assign J2END_CD_BEG3_input = {W2END0, S2END0, E2END0, N2END0};
  cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG3 (
      .A0 (J2END_CD_BEG3_input[0]),
      .A1 (J2END_CD_BEG3_input[1]),
      .A2 (J2END_CD_BEG3_input[2]),
      .A3 (J2END_CD_BEG3_input[3]),
      .S0 (ConfigBits[234+0]),
      .S0N(ConfigBits_N[234+0]),
      .S1 (ConfigBits[234+1]),
      .S1N(ConfigBits_N[234+1]),
      .X  (J2END_CD_BEG3)
  );

  // switch matrix multiplexer  J2END_EF_BEG0         MUX-4
  assign J2END_EF_BEG0_input = {W2END7, S2END7, E2END7, N2END7};
  cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG0 (
      .A0 (J2END_EF_BEG0_input[0]),
      .A1 (J2END_EF_BEG0_input[1]),
      .A2 (J2END_EF_BEG0_input[2]),
      .A3 (J2END_EF_BEG0_input[3]),
      .S0 (ConfigBits[236+0]),
      .S0N(ConfigBits_N[236+0]),
      .S1 (ConfigBits[236+1]),
      .S1N(ConfigBits_N[236+1]),
      .X  (J2END_EF_BEG0)
  );

  // switch matrix multiplexer  J2END_EF_BEG1         MUX-4
  assign J2END_EF_BEG1_input = {W2END3, S2END3, E2END3, N2END3};
  cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG1 (
      .A0 (J2END_EF_BEG1_input[0]),
      .A1 (J2END_EF_BEG1_input[1]),
      .A2 (J2END_EF_BEG1_input[2]),
      .A3 (J2END_EF_BEG1_input[3]),
      .S0 (ConfigBits[238+0]),
      .S0N(ConfigBits_N[238+0]),
      .S1 (ConfigBits[238+1]),
      .S1N(ConfigBits_N[238+1]),
      .X  (J2END_EF_BEG1)
  );

  // switch matrix multiplexer  J2END_EF_BEG2         MUX-4
  assign J2END_EF_BEG2_input = {W2END5, S2END5, E2END5, N2END5};
  cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG2 (
      .A0 (J2END_EF_BEG2_input[0]),
      .A1 (J2END_EF_BEG2_input[1]),
      .A2 (J2END_EF_BEG2_input[2]),
      .A3 (J2END_EF_BEG2_input[3]),
      .S0 (ConfigBits[240+0]),
      .S0N(ConfigBits_N[240+0]),
      .S1 (ConfigBits[240+1]),
      .S1N(ConfigBits_N[240+1]),
      .X  (J2END_EF_BEG2)
  );

  // switch matrix multiplexer  J2END_EF_BEG3         MUX-4
  assign J2END_EF_BEG3_input = {W2END1, S2END1, E2END1, N2END1};
  cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG3 (
      .A0 (J2END_EF_BEG3_input[0]),
      .A1 (J2END_EF_BEG3_input[1]),
      .A2 (J2END_EF_BEG3_input[2]),
      .A3 (J2END_EF_BEG3_input[3]),
      .S0 (ConfigBits[242+0]),
      .S0N(ConfigBits_N[242+0]),
      .S1 (ConfigBits[242+1]),
      .S1N(ConfigBits_N[242+1]),
      .X  (J2END_EF_BEG3)
  );

  // switch matrix multiplexer  J2END_GH_BEG0         MUX-4
  assign J2END_GH_BEG0_input = {W2END7, S2END7, E2END7, N2END7};
  cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG0 (
      .A0 (J2END_GH_BEG0_input[0]),
      .A1 (J2END_GH_BEG0_input[1]),
      .A2 (J2END_GH_BEG0_input[2]),
      .A3 (J2END_GH_BEG0_input[3]),
      .S0 (ConfigBits[244+0]),
      .S0N(ConfigBits_N[244+0]),
      .S1 (ConfigBits[244+1]),
      .S1N(ConfigBits_N[244+1]),
      .X  (J2END_GH_BEG0)
  );

  // switch matrix multiplexer  J2END_GH_BEG1         MUX-4
  assign J2END_GH_BEG1_input = {W2END3, S2END3, E2END3, N2END3};
  cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG1 (
      .A0 (J2END_GH_BEG1_input[0]),
      .A1 (J2END_GH_BEG1_input[1]),
      .A2 (J2END_GH_BEG1_input[2]),
      .A3 (J2END_GH_BEG1_input[3]),
      .S0 (ConfigBits[246+0]),
      .S0N(ConfigBits_N[246+0]),
      .S1 (ConfigBits[246+1]),
      .S1N(ConfigBits_N[246+1]),
      .X  (J2END_GH_BEG1)
  );

  // switch matrix multiplexer  J2END_GH_BEG2         MUX-4
  assign J2END_GH_BEG2_input = {W2END5, S2END5, E2END5, N2END5};
  cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG2 (
      .A0 (J2END_GH_BEG2_input[0]),
      .A1 (J2END_GH_BEG2_input[1]),
      .A2 (J2END_GH_BEG2_input[2]),
      .A3 (J2END_GH_BEG2_input[3]),
      .S0 (ConfigBits[248+0]),
      .S0N(ConfigBits_N[248+0]),
      .S1 (ConfigBits[248+1]),
      .S1N(ConfigBits_N[248+1]),
      .X  (J2END_GH_BEG2)
  );

  // switch matrix multiplexer  J2END_GH_BEG3         MUX-4
  assign J2END_GH_BEG3_input = {W2END1, S2END1, E2END1, N2END1};
  cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG3 (
      .A0 (J2END_GH_BEG3_input[0]),
      .A1 (J2END_GH_BEG3_input[1]),
      .A2 (J2END_GH_BEG3_input[2]),
      .A3 (J2END_GH_BEG3_input[3]),
      .S0 (ConfigBits[250+0]),
      .S0N(ConfigBits_N[250+0]),
      .S1 (ConfigBits[250+1]),
      .S1N(ConfigBits_N[250+1]),
      .X  (J2END_GH_BEG3)
  );

  // switch matrix multiplexer  JN2BEG0         MUX-16
  assign JN2BEG0_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    W6END1,
    W2END1,
    S2END1,
    E6END1,
    EE4END0,
    E2END1,
    E1END3,
    N4END1,
    N2END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG0 (
      .A0 (JN2BEG0_input[0]),
      .A1 (JN2BEG0_input[1]),
      .A2 (JN2BEG0_input[2]),
      .A3 (JN2BEG0_input[3]),
      .A4 (JN2BEG0_input[4]),
      .A5 (JN2BEG0_input[5]),
      .A6 (JN2BEG0_input[6]),
      .A7 (JN2BEG0_input[7]),
      .A8 (JN2BEG0_input[8]),
      .A9 (JN2BEG0_input[9]),
      .A10(JN2BEG0_input[10]),
      .A11(JN2BEG0_input[11]),
      .A12(JN2BEG0_input[12]),
      .A13(JN2BEG0_input[13]),
      .A14(JN2BEG0_input[14]),
      .A15(JN2BEG0_input[15]),
      .S0 (ConfigBits[252+0]),
      .S0N(ConfigBits_N[252+0]),
      .S1 (ConfigBits[252+1]),
      .S1N(ConfigBits_N[252+1]),
      .S2 (ConfigBits[252+2]),
      .S2N(ConfigBits_N[252+2]),
      .S3 (ConfigBits[252+3]),
      .S3N(ConfigBits_N[252+3]),
      .X  (JN2BEG0)
  );

  // switch matrix multiplexer  JN2BEG1         MUX-16
  assign JN2BEG1_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD0,
    W6END0,
    W2END2,
    S2END2,
    E6END0,
    EE4END1,
    E2END2,
    E1END0,
    N4END2,
    N2END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG1 (
      .A0 (JN2BEG1_input[0]),
      .A1 (JN2BEG1_input[1]),
      .A2 (JN2BEG1_input[2]),
      .A3 (JN2BEG1_input[3]),
      .A4 (JN2BEG1_input[4]),
      .A5 (JN2BEG1_input[5]),
      .A6 (JN2BEG1_input[6]),
      .A7 (JN2BEG1_input[7]),
      .A8 (JN2BEG1_input[8]),
      .A9 (JN2BEG1_input[9]),
      .A10(JN2BEG1_input[10]),
      .A11(JN2BEG1_input[11]),
      .A12(JN2BEG1_input[12]),
      .A13(JN2BEG1_input[13]),
      .A14(JN2BEG1_input[14]),
      .A15(JN2BEG1_input[15]),
      .S0 (ConfigBits[256+0]),
      .S0N(ConfigBits_N[256+0]),
      .S1 (ConfigBits[256+1]),
      .S1N(ConfigBits_N[256+1]),
      .S2 (ConfigBits[256+2]),
      .S2N(ConfigBits_N[256+2]),
      .S3 (ConfigBits[256+3]),
      .S3N(ConfigBits_N[256+3]),
      .X  (JN2BEG1)
  );

  // switch matrix multiplexer  JN2BEG2         MUX-16
  assign JN2BEG2_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD1,
    AD0,
    W6END1,
    WW4END2,
    W2END3,
    S2END3,
    E6END1,
    E2END3,
    E1END1,
    N4END3,
    N2END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG2 (
      .A0 (JN2BEG2_input[0]),
      .A1 (JN2BEG2_input[1]),
      .A2 (JN2BEG2_input[2]),
      .A3 (JN2BEG2_input[3]),
      .A4 (JN2BEG2_input[4]),
      .A5 (JN2BEG2_input[5]),
      .A6 (JN2BEG2_input[6]),
      .A7 (JN2BEG2_input[7]),
      .A8 (JN2BEG2_input[8]),
      .A9 (JN2BEG2_input[9]),
      .A10(JN2BEG2_input[10]),
      .A11(JN2BEG2_input[11]),
      .A12(JN2BEG2_input[12]),
      .A13(JN2BEG2_input[13]),
      .A14(JN2BEG2_input[14]),
      .A15(JN2BEG2_input[15]),
      .S0 (ConfigBits[260+0]),
      .S0N(ConfigBits_N[260+0]),
      .S1 (ConfigBits[260+1]),
      .S1N(ConfigBits_N[260+1]),
      .S2 (ConfigBits[260+2]),
      .S2N(ConfigBits_N[260+2]),
      .S3 (ConfigBits[260+3]),
      .S3N(ConfigBits_N[260+3]),
      .X  (JN2BEG2)
  );

  // switch matrix multiplexer  JN2BEG3         MUX-16
  assign JN2BEG3_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD2,
    AD1,
    AD0,
    W6END0,
    WW4END3,
    W2END4,
    S2END4,
    E6END0,
    E2END4,
    E1END2,
    N4END0,
    N2END4
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG3 (
      .A0 (JN2BEG3_input[0]),
      .A1 (JN2BEG3_input[1]),
      .A2 (JN2BEG3_input[2]),
      .A3 (JN2BEG3_input[3]),
      .A4 (JN2BEG3_input[4]),
      .A5 (JN2BEG3_input[5]),
      .A6 (JN2BEG3_input[6]),
      .A7 (JN2BEG3_input[7]),
      .A8 (JN2BEG3_input[8]),
      .A9 (JN2BEG3_input[9]),
      .A10(JN2BEG3_input[10]),
      .A11(JN2BEG3_input[11]),
      .A12(JN2BEG3_input[12]),
      .A13(JN2BEG3_input[13]),
      .A14(JN2BEG3_input[14]),
      .A15(JN2BEG3_input[15]),
      .S0 (ConfigBits[264+0]),
      .S0N(ConfigBits_N[264+0]),
      .S1 (ConfigBits[264+1]),
      .S1N(ConfigBits_N[264+1]),
      .S2 (ConfigBits[264+2]),
      .S2N(ConfigBits_N[264+2]),
      .S3 (ConfigBits[264+3]),
      .S3N(ConfigBits_N[264+3]),
      .X  (JN2BEG3)
  );

  // switch matrix multiplexer  JN2BEG4         MUX-16
  assign JN2BEG4_input = {
    BD3,
    BD2,
    BD1,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    W1END1,
    S2END5,
    S1END1,
    E2END5,
    E1END1,
    NN4END3,
    N2END5,
    N1END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG4 (
      .A0 (JN2BEG4_input[0]),
      .A1 (JN2BEG4_input[1]),
      .A2 (JN2BEG4_input[2]),
      .A3 (JN2BEG4_input[3]),
      .A4 (JN2BEG4_input[4]),
      .A5 (JN2BEG4_input[5]),
      .A6 (JN2BEG4_input[6]),
      .A7 (JN2BEG4_input[7]),
      .A8 (JN2BEG4_input[8]),
      .A9 (JN2BEG4_input[9]),
      .A10(JN2BEG4_input[10]),
      .A11(JN2BEG4_input[11]),
      .A12(JN2BEG4_input[12]),
      .A13(JN2BEG4_input[13]),
      .A14(JN2BEG4_input[14]),
      .A15(JN2BEG4_input[15]),
      .S0 (ConfigBits[268+0]),
      .S0N(ConfigBits_N[268+0]),
      .S1 (ConfigBits[268+1]),
      .S1N(ConfigBits_N[268+1]),
      .S2 (ConfigBits[268+2]),
      .S2N(ConfigBits_N[268+2]),
      .S3 (ConfigBits[268+3]),
      .S3N(ConfigBits_N[268+3]),
      .X  (JN2BEG4)
  );

  // switch matrix multiplexer  JN2BEG5         MUX-16
  assign JN2BEG5_input = {
    BD3,
    BD2,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    W1END0,
    S2END6,
    S1END2,
    E2END6,
    E1END2,
    NN4END2,
    N2END6,
    N1END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG5 (
      .A0 (JN2BEG5_input[0]),
      .A1 (JN2BEG5_input[1]),
      .A2 (JN2BEG5_input[2]),
      .A3 (JN2BEG5_input[3]),
      .A4 (JN2BEG5_input[4]),
      .A5 (JN2BEG5_input[5]),
      .A6 (JN2BEG5_input[6]),
      .A7 (JN2BEG5_input[7]),
      .A8 (JN2BEG5_input[8]),
      .A9 (JN2BEG5_input[9]),
      .A10(JN2BEG5_input[10]),
      .A11(JN2BEG5_input[11]),
      .A12(JN2BEG5_input[12]),
      .A13(JN2BEG5_input[13]),
      .A14(JN2BEG5_input[14]),
      .A15(JN2BEG5_input[15]),
      .S0 (ConfigBits[272+0]),
      .S0N(ConfigBits_N[272+0]),
      .S1 (ConfigBits[272+1]),
      .S1N(ConfigBits_N[272+1]),
      .S2 (ConfigBits[272+2]),
      .S2N(ConfigBits_N[272+2]),
      .S3 (ConfigBits[272+3]),
      .S3N(ConfigBits_N[272+3]),
      .X  (JN2BEG5)
  );

  // switch matrix multiplexer  JN2BEG6         MUX-16
  assign JN2BEG6_input = {
    BD3,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    W1END1,
    S2END7,
    S1END3,
    E2END7,
    E1END3,
    NN4END1,
    N2END7,
    N1END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG6 (
      .A0 (JN2BEG6_input[0]),
      .A1 (JN2BEG6_input[1]),
      .A2 (JN2BEG6_input[2]),
      .A3 (JN2BEG6_input[3]),
      .A4 (JN2BEG6_input[4]),
      .A5 (JN2BEG6_input[5]),
      .A6 (JN2BEG6_input[6]),
      .A7 (JN2BEG6_input[7]),
      .A8 (JN2BEG6_input[8]),
      .A9 (JN2BEG6_input[9]),
      .A10(JN2BEG6_input[10]),
      .A11(JN2BEG6_input[11]),
      .A12(JN2BEG6_input[12]),
      .A13(JN2BEG6_input[13]),
      .A14(JN2BEG6_input[14]),
      .A15(JN2BEG6_input[15]),
      .S0 (ConfigBits[276+0]),
      .S0N(ConfigBits_N[276+0]),
      .S1 (ConfigBits[276+1]),
      .S1N(ConfigBits_N[276+1]),
      .S2 (ConfigBits[276+2]),
      .S2N(ConfigBits_N[276+2]),
      .S3 (ConfigBits[276+3]),
      .S3N(ConfigBits_N[276+3]),
      .X  (JN2BEG6)
  );

  // switch matrix multiplexer  JN2BEG7         MUX-16
  assign JN2BEG7_input = {
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    W1END0,
    S2END0,
    S1END0,
    E2END0,
    E1END0,
    NN4END0,
    N2END0,
    N1END0
  };
  cus_mux161_buf inst_cus_mux161_buf_JN2BEG7 (
      .A0 (JN2BEG7_input[0]),
      .A1 (JN2BEG7_input[1]),
      .A2 (JN2BEG7_input[2]),
      .A3 (JN2BEG7_input[3]),
      .A4 (JN2BEG7_input[4]),
      .A5 (JN2BEG7_input[5]),
      .A6 (JN2BEG7_input[6]),
      .A7 (JN2BEG7_input[7]),
      .A8 (JN2BEG7_input[8]),
      .A9 (JN2BEG7_input[9]),
      .A10(JN2BEG7_input[10]),
      .A11(JN2BEG7_input[11]),
      .A12(JN2BEG7_input[12]),
      .A13(JN2BEG7_input[13]),
      .A14(JN2BEG7_input[14]),
      .A15(JN2BEG7_input[15]),
      .S0 (ConfigBits[280+0]),
      .S0N(ConfigBits_N[280+0]),
      .S1 (ConfigBits[280+1]),
      .S1N(ConfigBits_N[280+1]),
      .S2 (ConfigBits[280+2]),
      .S2N(ConfigBits_N[280+2]),
      .S3 (ConfigBits[280+3]),
      .S3N(ConfigBits_N[280+3]),
      .X  (JN2BEG7)
  );

  // switch matrix multiplexer  JE2BEG0         MUX-16
  assign JE2BEG0_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    W6END1,
    W2END1,
    S2END1,
    E6END1,
    E2END1,
    NN4END0,
    N4END1,
    N2END1,
    N1END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG0 (
      .A0 (JE2BEG0_input[0]),
      .A1 (JE2BEG0_input[1]),
      .A2 (JE2BEG0_input[2]),
      .A3 (JE2BEG0_input[3]),
      .A4 (JE2BEG0_input[4]),
      .A5 (JE2BEG0_input[5]),
      .A6 (JE2BEG0_input[6]),
      .A7 (JE2BEG0_input[7]),
      .A8 (JE2BEG0_input[8]),
      .A9 (JE2BEG0_input[9]),
      .A10(JE2BEG0_input[10]),
      .A11(JE2BEG0_input[11]),
      .A12(JE2BEG0_input[12]),
      .A13(JE2BEG0_input[13]),
      .A14(JE2BEG0_input[14]),
      .A15(JE2BEG0_input[15]),
      .S0 (ConfigBits[284+0]),
      .S0N(ConfigBits_N[284+0]),
      .S1 (ConfigBits[284+1]),
      .S1N(ConfigBits_N[284+1]),
      .S2 (ConfigBits[284+2]),
      .S2N(ConfigBits_N[284+2]),
      .S3 (ConfigBits[284+3]),
      .S3N(ConfigBits_N[284+3]),
      .X  (JE2BEG0)
  );

  // switch matrix multiplexer  JE2BEG1         MUX-16
  assign JE2BEG1_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD0,
    W6END0,
    W2END2,
    S2END2,
    E6END0,
    E2END2,
    NN4END1,
    N4END2,
    N2END2,
    N1END0
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG1 (
      .A0 (JE2BEG1_input[0]),
      .A1 (JE2BEG1_input[1]),
      .A2 (JE2BEG1_input[2]),
      .A3 (JE2BEG1_input[3]),
      .A4 (JE2BEG1_input[4]),
      .A5 (JE2BEG1_input[5]),
      .A6 (JE2BEG1_input[6]),
      .A7 (JE2BEG1_input[7]),
      .A8 (JE2BEG1_input[8]),
      .A9 (JE2BEG1_input[9]),
      .A10(JE2BEG1_input[10]),
      .A11(JE2BEG1_input[11]),
      .A12(JE2BEG1_input[12]),
      .A13(JE2BEG1_input[13]),
      .A14(JE2BEG1_input[14]),
      .A15(JE2BEG1_input[15]),
      .S0 (ConfigBits[288+0]),
      .S0N(ConfigBits_N[288+0]),
      .S1 (ConfigBits[288+1]),
      .S1N(ConfigBits_N[288+1]),
      .S2 (ConfigBits[288+2]),
      .S2N(ConfigBits_N[288+2]),
      .S3 (ConfigBits[288+3]),
      .S3N(ConfigBits_N[288+3]),
      .X  (JE2BEG1)
  );

  // switch matrix multiplexer  JE2BEG2         MUX-16
  assign JE2BEG2_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD1,
    AD0,
    W6END1,
    W2END3,
    SS4END2,
    S2END3,
    E6END1,
    E2END3,
    N4END3,
    N2END3,
    N1END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG2 (
      .A0 (JE2BEG2_input[0]),
      .A1 (JE2BEG2_input[1]),
      .A2 (JE2BEG2_input[2]),
      .A3 (JE2BEG2_input[3]),
      .A4 (JE2BEG2_input[4]),
      .A5 (JE2BEG2_input[5]),
      .A6 (JE2BEG2_input[6]),
      .A7 (JE2BEG2_input[7]),
      .A8 (JE2BEG2_input[8]),
      .A9 (JE2BEG2_input[9]),
      .A10(JE2BEG2_input[10]),
      .A11(JE2BEG2_input[11]),
      .A12(JE2BEG2_input[12]),
      .A13(JE2BEG2_input[13]),
      .A14(JE2BEG2_input[14]),
      .A15(JE2BEG2_input[15]),
      .S0 (ConfigBits[292+0]),
      .S0N(ConfigBits_N[292+0]),
      .S1 (ConfigBits[292+1]),
      .S1N(ConfigBits_N[292+1]),
      .S2 (ConfigBits[292+2]),
      .S2N(ConfigBits_N[292+2]),
      .S3 (ConfigBits[292+3]),
      .S3N(ConfigBits_N[292+3]),
      .X  (JE2BEG2)
  );

  // switch matrix multiplexer  JE2BEG3         MUX-16
  assign JE2BEG3_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD2,
    AD1,
    AD0,
    W6END0,
    W2END4,
    SS4END3,
    S2END4,
    E6END0,
    E2END4,
    N4END0,
    N2END4,
    N1END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG3 (
      .A0 (JE2BEG3_input[0]),
      .A1 (JE2BEG3_input[1]),
      .A2 (JE2BEG3_input[2]),
      .A3 (JE2BEG3_input[3]),
      .A4 (JE2BEG3_input[4]),
      .A5 (JE2BEG3_input[5]),
      .A6 (JE2BEG3_input[6]),
      .A7 (JE2BEG3_input[7]),
      .A8 (JE2BEG3_input[8]),
      .A9 (JE2BEG3_input[9]),
      .A10(JE2BEG3_input[10]),
      .A11(JE2BEG3_input[11]),
      .A12(JE2BEG3_input[12]),
      .A13(JE2BEG3_input[13]),
      .A14(JE2BEG3_input[14]),
      .A15(JE2BEG3_input[15]),
      .S0 (ConfigBits[296+0]),
      .S0N(ConfigBits_N[296+0]),
      .S1 (ConfigBits[296+1]),
      .S1N(ConfigBits_N[296+1]),
      .S2 (ConfigBits[296+2]),
      .S2N(ConfigBits_N[296+2]),
      .S3 (ConfigBits[296+3]),
      .S3N(ConfigBits_N[296+3]),
      .X  (JE2BEG3)
  );

  // switch matrix multiplexer  JE2BEG4         MUX-16
  assign JE2BEG4_input = {
    BD3,
    BD2,
    BD1,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END1,
    S2END5,
    S1END3,
    S1END1,
    EE4END3,
    E2END5,
    E1END1,
    N2END5,
    N1END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG4 (
      .A0 (JE2BEG4_input[0]),
      .A1 (JE2BEG4_input[1]),
      .A2 (JE2BEG4_input[2]),
      .A3 (JE2BEG4_input[3]),
      .A4 (JE2BEG4_input[4]),
      .A5 (JE2BEG4_input[5]),
      .A6 (JE2BEG4_input[6]),
      .A7 (JE2BEG4_input[7]),
      .A8 (JE2BEG4_input[8]),
      .A9 (JE2BEG4_input[9]),
      .A10(JE2BEG4_input[10]),
      .A11(JE2BEG4_input[11]),
      .A12(JE2BEG4_input[12]),
      .A13(JE2BEG4_input[13]),
      .A14(JE2BEG4_input[14]),
      .A15(JE2BEG4_input[15]),
      .S0 (ConfigBits[300+0]),
      .S0N(ConfigBits_N[300+0]),
      .S1 (ConfigBits[300+1]),
      .S1N(ConfigBits_N[300+1]),
      .S2 (ConfigBits[300+2]),
      .S2N(ConfigBits_N[300+2]),
      .S3 (ConfigBits[300+3]),
      .S3N(ConfigBits_N[300+3]),
      .X  (JE2BEG4)
  );

  // switch matrix multiplexer  JE2BEG5         MUX-16
  assign JE2BEG5_input = {
    BD3,
    BD2,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    S2END6,
    S1END2,
    S1END0,
    EE4END2,
    E2END6,
    E1END2,
    N2END6,
    N1END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG5 (
      .A0 (JE2BEG5_input[0]),
      .A1 (JE2BEG5_input[1]),
      .A2 (JE2BEG5_input[2]),
      .A3 (JE2BEG5_input[3]),
      .A4 (JE2BEG5_input[4]),
      .A5 (JE2BEG5_input[5]),
      .A6 (JE2BEG5_input[6]),
      .A7 (JE2BEG5_input[7]),
      .A8 (JE2BEG5_input[8]),
      .A9 (JE2BEG5_input[9]),
      .A10(JE2BEG5_input[10]),
      .A11(JE2BEG5_input[11]),
      .A12(JE2BEG5_input[12]),
      .A13(JE2BEG5_input[13]),
      .A14(JE2BEG5_input[14]),
      .A15(JE2BEG5_input[15]),
      .S0 (ConfigBits[304+0]),
      .S0N(ConfigBits_N[304+0]),
      .S1 (ConfigBits[304+1]),
      .S1N(ConfigBits_N[304+1]),
      .S2 (ConfigBits[304+2]),
      .S2N(ConfigBits_N[304+2]),
      .S3 (ConfigBits[304+3]),
      .S3N(ConfigBits_N[304+3]),
      .X  (JE2BEG5)
  );

  // switch matrix multiplexer  JE2BEG6         MUX-16
  assign JE2BEG6_input = {
    BD3,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    S2END7,
    S1END3,
    S1END1,
    EE4END1,
    E2END7,
    E1END3,
    N2END7,
    N1END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG6 (
      .A0 (JE2BEG6_input[0]),
      .A1 (JE2BEG6_input[1]),
      .A2 (JE2BEG6_input[2]),
      .A3 (JE2BEG6_input[3]),
      .A4 (JE2BEG6_input[4]),
      .A5 (JE2BEG6_input[5]),
      .A6 (JE2BEG6_input[6]),
      .A7 (JE2BEG6_input[7]),
      .A8 (JE2BEG6_input[8]),
      .A9 (JE2BEG6_input[9]),
      .A10(JE2BEG6_input[10]),
      .A11(JE2BEG6_input[11]),
      .A12(JE2BEG6_input[12]),
      .A13(JE2BEG6_input[13]),
      .A14(JE2BEG6_input[14]),
      .A15(JE2BEG6_input[15]),
      .S0 (ConfigBits[308+0]),
      .S0N(ConfigBits_N[308+0]),
      .S1 (ConfigBits[308+1]),
      .S1N(ConfigBits_N[308+1]),
      .S2 (ConfigBits[308+2]),
      .S2N(ConfigBits_N[308+2]),
      .S3 (ConfigBits[308+3]),
      .S3N(ConfigBits_N[308+3]),
      .X  (JE2BEG6)
  );

  // switch matrix multiplexer  JE2BEG7         MUX-16
  assign JE2BEG7_input = {
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END0,
    S2END0,
    S1END2,
    S1END0,
    EE4END0,
    E2END0,
    E1END0,
    N2END0,
    N1END0
  };
  cus_mux161_buf inst_cus_mux161_buf_JE2BEG7 (
      .A0 (JE2BEG7_input[0]),
      .A1 (JE2BEG7_input[1]),
      .A2 (JE2BEG7_input[2]),
      .A3 (JE2BEG7_input[3]),
      .A4 (JE2BEG7_input[4]),
      .A5 (JE2BEG7_input[5]),
      .A6 (JE2BEG7_input[6]),
      .A7 (JE2BEG7_input[7]),
      .A8 (JE2BEG7_input[8]),
      .A9 (JE2BEG7_input[9]),
      .A10(JE2BEG7_input[10]),
      .A11(JE2BEG7_input[11]),
      .A12(JE2BEG7_input[12]),
      .A13(JE2BEG7_input[13]),
      .A14(JE2BEG7_input[14]),
      .A15(JE2BEG7_input[15]),
      .S0 (ConfigBits[312+0]),
      .S0N(ConfigBits_N[312+0]),
      .S1 (ConfigBits[312+1]),
      .S1N(ConfigBits_N[312+1]),
      .S2 (ConfigBits[312+2]),
      .S2N(ConfigBits_N[312+2]),
      .S3 (ConfigBits[312+3]),
      .S3N(ConfigBits_N[312+3]),
      .X  (JE2BEG7)
  );

  // switch matrix multiplexer  JS2BEG0         MUX-16
  assign JS2BEG0_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    W6END1,
    WW4END0,
    W2END1,
    S4END1,
    S2END1,
    E6END1,
    E2END1,
    E1END3,
    N2END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG0 (
      .A0 (JS2BEG0_input[0]),
      .A1 (JS2BEG0_input[1]),
      .A2 (JS2BEG0_input[2]),
      .A3 (JS2BEG0_input[3]),
      .A4 (JS2BEG0_input[4]),
      .A5 (JS2BEG0_input[5]),
      .A6 (JS2BEG0_input[6]),
      .A7 (JS2BEG0_input[7]),
      .A8 (JS2BEG0_input[8]),
      .A9 (JS2BEG0_input[9]),
      .A10(JS2BEG0_input[10]),
      .A11(JS2BEG0_input[11]),
      .A12(JS2BEG0_input[12]),
      .A13(JS2BEG0_input[13]),
      .A14(JS2BEG0_input[14]),
      .A15(JS2BEG0_input[15]),
      .S0 (ConfigBits[316+0]),
      .S0N(ConfigBits_N[316+0]),
      .S1 (ConfigBits[316+1]),
      .S1N(ConfigBits_N[316+1]),
      .S2 (ConfigBits[316+2]),
      .S2N(ConfigBits_N[316+2]),
      .S3 (ConfigBits[316+3]),
      .S3N(ConfigBits_N[316+3]),
      .X  (JS2BEG0)
  );

  // switch matrix multiplexer  JS2BEG1         MUX-16
  assign JS2BEG1_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD0,
    W6END0,
    WW4END1,
    W2END2,
    S4END2,
    S2END2,
    E6END0,
    E2END2,
    E1END0,
    N2END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG1 (
      .A0 (JS2BEG1_input[0]),
      .A1 (JS2BEG1_input[1]),
      .A2 (JS2BEG1_input[2]),
      .A3 (JS2BEG1_input[3]),
      .A4 (JS2BEG1_input[4]),
      .A5 (JS2BEG1_input[5]),
      .A6 (JS2BEG1_input[6]),
      .A7 (JS2BEG1_input[7]),
      .A8 (JS2BEG1_input[8]),
      .A9 (JS2BEG1_input[9]),
      .A10(JS2BEG1_input[10]),
      .A11(JS2BEG1_input[11]),
      .A12(JS2BEG1_input[12]),
      .A13(JS2BEG1_input[13]),
      .A14(JS2BEG1_input[14]),
      .A15(JS2BEG1_input[15]),
      .S0 (ConfigBits[320+0]),
      .S0N(ConfigBits_N[320+0]),
      .S1 (ConfigBits[320+1]),
      .S1N(ConfigBits_N[320+1]),
      .S2 (ConfigBits[320+2]),
      .S2N(ConfigBits_N[320+2]),
      .S3 (ConfigBits[320+3]),
      .S3N(ConfigBits_N[320+3]),
      .X  (JS2BEG1)
  );

  // switch matrix multiplexer  JS2BEG2         MUX-16
  assign JS2BEG2_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD1,
    AD0,
    W6END1,
    W2END3,
    S4END3,
    S2END3,
    E6END1,
    EE4END2,
    E2END3,
    E1END1,
    N2END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG2 (
      .A0 (JS2BEG2_input[0]),
      .A1 (JS2BEG2_input[1]),
      .A2 (JS2BEG2_input[2]),
      .A3 (JS2BEG2_input[3]),
      .A4 (JS2BEG2_input[4]),
      .A5 (JS2BEG2_input[5]),
      .A6 (JS2BEG2_input[6]),
      .A7 (JS2BEG2_input[7]),
      .A8 (JS2BEG2_input[8]),
      .A9 (JS2BEG2_input[9]),
      .A10(JS2BEG2_input[10]),
      .A11(JS2BEG2_input[11]),
      .A12(JS2BEG2_input[12]),
      .A13(JS2BEG2_input[13]),
      .A14(JS2BEG2_input[14]),
      .A15(JS2BEG2_input[15]),
      .S0 (ConfigBits[324+0]),
      .S0N(ConfigBits_N[324+0]),
      .S1 (ConfigBits[324+1]),
      .S1N(ConfigBits_N[324+1]),
      .S2 (ConfigBits[324+2]),
      .S2N(ConfigBits_N[324+2]),
      .S3 (ConfigBits[324+3]),
      .S3N(ConfigBits_N[324+3]),
      .X  (JS2BEG2)
  );

  // switch matrix multiplexer  JS2BEG3         MUX-16
  assign JS2BEG3_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD2,
    AD1,
    AD0,
    W6END0,
    W2END4,
    S4END0,
    S2END4,
    E6END0,
    EE4END3,
    E2END4,
    E1END2,
    N2END4
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG3 (
      .A0 (JS2BEG3_input[0]),
      .A1 (JS2BEG3_input[1]),
      .A2 (JS2BEG3_input[2]),
      .A3 (JS2BEG3_input[3]),
      .A4 (JS2BEG3_input[4]),
      .A5 (JS2BEG3_input[5]),
      .A6 (JS2BEG3_input[6]),
      .A7 (JS2BEG3_input[7]),
      .A8 (JS2BEG3_input[8]),
      .A9 (JS2BEG3_input[9]),
      .A10(JS2BEG3_input[10]),
      .A11(JS2BEG3_input[11]),
      .A12(JS2BEG3_input[12]),
      .A13(JS2BEG3_input[13]),
      .A14(JS2BEG3_input[14]),
      .A15(JS2BEG3_input[15]),
      .S0 (ConfigBits[328+0]),
      .S0N(ConfigBits_N[328+0]),
      .S1 (ConfigBits[328+1]),
      .S1N(ConfigBits_N[328+1]),
      .S2 (ConfigBits[328+2]),
      .S2N(ConfigBits_N[328+2]),
      .S3 (ConfigBits[328+3]),
      .S3N(ConfigBits_N[328+3]),
      .X  (JS2BEG3)
  );

  // switch matrix multiplexer  JS2BEG4         MUX-16
  assign JS2BEG4_input = {
    BD3,
    BD2,
    BD1,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    W1END1,
    SS4END3,
    S2END5,
    S1END1,
    E2END5,
    E1END1,
    N2END5,
    N1END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG4 (
      .A0 (JS2BEG4_input[0]),
      .A1 (JS2BEG4_input[1]),
      .A2 (JS2BEG4_input[2]),
      .A3 (JS2BEG4_input[3]),
      .A4 (JS2BEG4_input[4]),
      .A5 (JS2BEG4_input[5]),
      .A6 (JS2BEG4_input[6]),
      .A7 (JS2BEG4_input[7]),
      .A8 (JS2BEG4_input[8]),
      .A9 (JS2BEG4_input[9]),
      .A10(JS2BEG4_input[10]),
      .A11(JS2BEG4_input[11]),
      .A12(JS2BEG4_input[12]),
      .A13(JS2BEG4_input[13]),
      .A14(JS2BEG4_input[14]),
      .A15(JS2BEG4_input[15]),
      .S0 (ConfigBits[332+0]),
      .S0N(ConfigBits_N[332+0]),
      .S1 (ConfigBits[332+1]),
      .S1N(ConfigBits_N[332+1]),
      .S2 (ConfigBits[332+2]),
      .S2N(ConfigBits_N[332+2]),
      .S3 (ConfigBits[332+3]),
      .S3N(ConfigBits_N[332+3]),
      .X  (JS2BEG4)
  );

  // switch matrix multiplexer  JS2BEG5         MUX-16
  assign JS2BEG5_input = {
    BD3,
    BD2,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    W1END0,
    SS4END2,
    S2END6,
    S1END2,
    E2END6,
    E1END2,
    N2END6,
    N1END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG5 (
      .A0 (JS2BEG5_input[0]),
      .A1 (JS2BEG5_input[1]),
      .A2 (JS2BEG5_input[2]),
      .A3 (JS2BEG5_input[3]),
      .A4 (JS2BEG5_input[4]),
      .A5 (JS2BEG5_input[5]),
      .A6 (JS2BEG5_input[6]),
      .A7 (JS2BEG5_input[7]),
      .A8 (JS2BEG5_input[8]),
      .A9 (JS2BEG5_input[9]),
      .A10(JS2BEG5_input[10]),
      .A11(JS2BEG5_input[11]),
      .A12(JS2BEG5_input[12]),
      .A13(JS2BEG5_input[13]),
      .A14(JS2BEG5_input[14]),
      .A15(JS2BEG5_input[15]),
      .S0 (ConfigBits[336+0]),
      .S0N(ConfigBits_N[336+0]),
      .S1 (ConfigBits[336+1]),
      .S1N(ConfigBits_N[336+1]),
      .S2 (ConfigBits[336+2]),
      .S2N(ConfigBits_N[336+2]),
      .S3 (ConfigBits[336+3]),
      .S3N(ConfigBits_N[336+3]),
      .X  (JS2BEG5)
  );

  // switch matrix multiplexer  JS2BEG6         MUX-16
  assign JS2BEG6_input = {
    BD3,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END3,
    W1END1,
    SS4END1,
    S2END7,
    S1END3,
    E2END7,
    E1END3,
    N2END7,
    N1END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG6 (
      .A0 (JS2BEG6_input[0]),
      .A1 (JS2BEG6_input[1]),
      .A2 (JS2BEG6_input[2]),
      .A3 (JS2BEG6_input[3]),
      .A4 (JS2BEG6_input[4]),
      .A5 (JS2BEG6_input[5]),
      .A6 (JS2BEG6_input[6]),
      .A7 (JS2BEG6_input[7]),
      .A8 (JS2BEG6_input[8]),
      .A9 (JS2BEG6_input[9]),
      .A10(JS2BEG6_input[10]),
      .A11(JS2BEG6_input[11]),
      .A12(JS2BEG6_input[12]),
      .A13(JS2BEG6_input[13]),
      .A14(JS2BEG6_input[14]),
      .A15(JS2BEG6_input[15]),
      .S0 (ConfigBits[340+0]),
      .S0N(ConfigBits_N[340+0]),
      .S1 (ConfigBits[340+1]),
      .S1N(ConfigBits_N[340+1]),
      .S2 (ConfigBits[340+2]),
      .S2N(ConfigBits_N[340+2]),
      .S3 (ConfigBits[340+3]),
      .S3N(ConfigBits_N[340+3]),
      .X  (JS2BEG6)
  );

  // switch matrix multiplexer  JS2BEG7         MUX-16
  assign JS2BEG7_input = {
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    W1END2,
    W1END0,
    SS4END0,
    S2END0,
    S1END0,
    E2END0,
    E1END0,
    N2END0,
    N1END0
  };
  cus_mux161_buf inst_cus_mux161_buf_JS2BEG7 (
      .A0 (JS2BEG7_input[0]),
      .A1 (JS2BEG7_input[1]),
      .A2 (JS2BEG7_input[2]),
      .A3 (JS2BEG7_input[3]),
      .A4 (JS2BEG7_input[4]),
      .A5 (JS2BEG7_input[5]),
      .A6 (JS2BEG7_input[6]),
      .A7 (JS2BEG7_input[7]),
      .A8 (JS2BEG7_input[8]),
      .A9 (JS2BEG7_input[9]),
      .A10(JS2BEG7_input[10]),
      .A11(JS2BEG7_input[11]),
      .A12(JS2BEG7_input[12]),
      .A13(JS2BEG7_input[13]),
      .A14(JS2BEG7_input[14]),
      .A15(JS2BEG7_input[15]),
      .S0 (ConfigBits[344+0]),
      .S0N(ConfigBits_N[344+0]),
      .S1 (ConfigBits[344+1]),
      .S1N(ConfigBits_N[344+1]),
      .S2 (ConfigBits[344+2]),
      .S2N(ConfigBits_N[344+2]),
      .S3 (ConfigBits[344+3]),
      .S3N(ConfigBits_N[344+3]),
      .X  (JS2BEG7)
  );

  // switch matrix multiplexer  JW2BEG0         MUX-16
  assign JW2BEG0_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    W6END1,
    W2END1,
    SS4END0,
    S4END1,
    S2END1,
    E6END1,
    E2END1,
    N2END1,
    N1END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG0 (
      .A0 (JW2BEG0_input[0]),
      .A1 (JW2BEG0_input[1]),
      .A2 (JW2BEG0_input[2]),
      .A3 (JW2BEG0_input[3]),
      .A4 (JW2BEG0_input[4]),
      .A5 (JW2BEG0_input[5]),
      .A6 (JW2BEG0_input[6]),
      .A7 (JW2BEG0_input[7]),
      .A8 (JW2BEG0_input[8]),
      .A9 (JW2BEG0_input[9]),
      .A10(JW2BEG0_input[10]),
      .A11(JW2BEG0_input[11]),
      .A12(JW2BEG0_input[12]),
      .A13(JW2BEG0_input[13]),
      .A14(JW2BEG0_input[14]),
      .A15(JW2BEG0_input[15]),
      .S0 (ConfigBits[348+0]),
      .S0N(ConfigBits_N[348+0]),
      .S1 (ConfigBits[348+1]),
      .S1N(ConfigBits_N[348+1]),
      .S2 (ConfigBits[348+2]),
      .S2N(ConfigBits_N[348+2]),
      .S3 (ConfigBits[348+3]),
      .S3N(ConfigBits_N[348+3]),
      .X  (JW2BEG0)
  );

  // switch matrix multiplexer  JW2BEG1         MUX-16
  assign JW2BEG1_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD0,
    W6END0,
    W2END2,
    SS4END1,
    S4END2,
    S2END2,
    E6END0,
    E2END2,
    N2END2,
    N1END0
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG1 (
      .A0 (JW2BEG1_input[0]),
      .A1 (JW2BEG1_input[1]),
      .A2 (JW2BEG1_input[2]),
      .A3 (JW2BEG1_input[3]),
      .A4 (JW2BEG1_input[4]),
      .A5 (JW2BEG1_input[5]),
      .A6 (JW2BEG1_input[6]),
      .A7 (JW2BEG1_input[7]),
      .A8 (JW2BEG1_input[8]),
      .A9 (JW2BEG1_input[9]),
      .A10(JW2BEG1_input[10]),
      .A11(JW2BEG1_input[11]),
      .A12(JW2BEG1_input[12]),
      .A13(JW2BEG1_input[13]),
      .A14(JW2BEG1_input[14]),
      .A15(JW2BEG1_input[15]),
      .S0 (ConfigBits[352+0]),
      .S0N(ConfigBits_N[352+0]),
      .S1 (ConfigBits[352+1]),
      .S1N(ConfigBits_N[352+1]),
      .S2 (ConfigBits[352+2]),
      .S2N(ConfigBits_N[352+2]),
      .S3 (ConfigBits[352+3]),
      .S3N(ConfigBits_N[352+3]),
      .X  (JW2BEG1)
  );

  // switch matrix multiplexer  JW2BEG2         MUX-16
  assign JW2BEG2_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD3,
    AD1,
    AD0,
    W6END1,
    W2END3,
    S4END3,
    S2END3,
    E6END1,
    E2END3,
    NN4END2,
    N2END3,
    N1END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG2 (
      .A0 (JW2BEG2_input[0]),
      .A1 (JW2BEG2_input[1]),
      .A2 (JW2BEG2_input[2]),
      .A3 (JW2BEG2_input[3]),
      .A4 (JW2BEG2_input[4]),
      .A5 (JW2BEG2_input[5]),
      .A6 (JW2BEG2_input[6]),
      .A7 (JW2BEG2_input[7]),
      .A8 (JW2BEG2_input[8]),
      .A9 (JW2BEG2_input[9]),
      .A10(JW2BEG2_input[10]),
      .A11(JW2BEG2_input[11]),
      .A12(JW2BEG2_input[12]),
      .A13(JW2BEG2_input[13]),
      .A14(JW2BEG2_input[14]),
      .A15(JW2BEG2_input[15]),
      .S0 (ConfigBits[356+0]),
      .S0N(ConfigBits_N[356+0]),
      .S1 (ConfigBits[356+1]),
      .S1N(ConfigBits_N[356+1]),
      .S2 (ConfigBits[356+2]),
      .S2N(ConfigBits_N[356+2]),
      .S3 (ConfigBits[356+3]),
      .S3N(ConfigBits_N[356+3]),
      .X  (JW2BEG2)
  );

  // switch matrix multiplexer  JW2BEG3         MUX-16
  assign JW2BEG3_input = {
    BD3,
    BD2,
    BD1,
    BD0,
    AD2,
    AD1,
    AD0,
    W6END0,
    W2END4,
    S4END0,
    S2END4,
    E6END0,
    E2END4,
    NN4END3,
    N2END4,
    N1END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG3 (
      .A0 (JW2BEG3_input[0]),
      .A1 (JW2BEG3_input[1]),
      .A2 (JW2BEG3_input[2]),
      .A3 (JW2BEG3_input[3]),
      .A4 (JW2BEG3_input[4]),
      .A5 (JW2BEG3_input[5]),
      .A6 (JW2BEG3_input[6]),
      .A7 (JW2BEG3_input[7]),
      .A8 (JW2BEG3_input[8]),
      .A9 (JW2BEG3_input[9]),
      .A10(JW2BEG3_input[10]),
      .A11(JW2BEG3_input[11]),
      .A12(JW2BEG3_input[12]),
      .A13(JW2BEG3_input[13]),
      .A14(JW2BEG3_input[14]),
      .A15(JW2BEG3_input[15]),
      .S0 (ConfigBits[360+0]),
      .S0N(ConfigBits_N[360+0]),
      .S1 (ConfigBits[360+1]),
      .S1N(ConfigBits_N[360+1]),
      .S2 (ConfigBits[360+2]),
      .S2N(ConfigBits_N[360+2]),
      .S3 (ConfigBits[360+3]),
      .S3N(ConfigBits_N[360+3]),
      .X  (JW2BEG3)
  );

  // switch matrix multiplexer  JW2BEG4         MUX-16
  assign JW2BEG4_input = {
    BD3,
    BD2,
    BD1,
    AD3,
    AD2,
    AD1,
    AD0,
    WW4END3,
    W1END1,
    S2END5,
    S1END3,
    S1END1,
    E2END5,
    E1END1,
    N2END5,
    N1END1
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG4 (
      .A0 (JW2BEG4_input[0]),
      .A1 (JW2BEG4_input[1]),
      .A2 (JW2BEG4_input[2]),
      .A3 (JW2BEG4_input[3]),
      .A4 (JW2BEG4_input[4]),
      .A5 (JW2BEG4_input[5]),
      .A6 (JW2BEG4_input[6]),
      .A7 (JW2BEG4_input[7]),
      .A8 (JW2BEG4_input[8]),
      .A9 (JW2BEG4_input[9]),
      .A10(JW2BEG4_input[10]),
      .A11(JW2BEG4_input[11]),
      .A12(JW2BEG4_input[12]),
      .A13(JW2BEG4_input[13]),
      .A14(JW2BEG4_input[14]),
      .A15(JW2BEG4_input[15]),
      .S0 (ConfigBits[364+0]),
      .S0N(ConfigBits_N[364+0]),
      .S1 (ConfigBits[364+1]),
      .S1N(ConfigBits_N[364+1]),
      .S2 (ConfigBits[364+2]),
      .S2N(ConfigBits_N[364+2]),
      .S3 (ConfigBits[364+3]),
      .S3N(ConfigBits_N[364+3]),
      .X  (JW2BEG4)
  );

  // switch matrix multiplexer  JW2BEG5         MUX-16
  assign JW2BEG5_input = {
    BD3,
    BD2,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    WW4END2,
    W1END2,
    S2END6,
    S1END2,
    S1END0,
    E2END6,
    E1END2,
    N2END6,
    N1END2
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG5 (
      .A0 (JW2BEG5_input[0]),
      .A1 (JW2BEG5_input[1]),
      .A2 (JW2BEG5_input[2]),
      .A3 (JW2BEG5_input[3]),
      .A4 (JW2BEG5_input[4]),
      .A5 (JW2BEG5_input[5]),
      .A6 (JW2BEG5_input[6]),
      .A7 (JW2BEG5_input[7]),
      .A8 (JW2BEG5_input[8]),
      .A9 (JW2BEG5_input[9]),
      .A10(JW2BEG5_input[10]),
      .A11(JW2BEG5_input[11]),
      .A12(JW2BEG5_input[12]),
      .A13(JW2BEG5_input[13]),
      .A14(JW2BEG5_input[14]),
      .A15(JW2BEG5_input[15]),
      .S0 (ConfigBits[368+0]),
      .S0N(ConfigBits_N[368+0]),
      .S1 (ConfigBits[368+1]),
      .S1N(ConfigBits_N[368+1]),
      .S2 (ConfigBits[368+2]),
      .S2N(ConfigBits_N[368+2]),
      .S3 (ConfigBits[368+3]),
      .S3N(ConfigBits_N[368+3]),
      .X  (JW2BEG5)
  );

  // switch matrix multiplexer  JW2BEG6         MUX-16
  assign JW2BEG6_input = {
    BD3,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    WW4END1,
    W1END3,
    S2END7,
    S1END3,
    S1END1,
    E2END7,
    E1END3,
    N2END7,
    N1END3
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG6 (
      .A0 (JW2BEG6_input[0]),
      .A1 (JW2BEG6_input[1]),
      .A2 (JW2BEG6_input[2]),
      .A3 (JW2BEG6_input[3]),
      .A4 (JW2BEG6_input[4]),
      .A5 (JW2BEG6_input[5]),
      .A6 (JW2BEG6_input[6]),
      .A7 (JW2BEG6_input[7]),
      .A8 (JW2BEG6_input[8]),
      .A9 (JW2BEG6_input[9]),
      .A10(JW2BEG6_input[10]),
      .A11(JW2BEG6_input[11]),
      .A12(JW2BEG6_input[12]),
      .A13(JW2BEG6_input[13]),
      .A14(JW2BEG6_input[14]),
      .A15(JW2BEG6_input[15]),
      .S0 (ConfigBits[372+0]),
      .S0N(ConfigBits_N[372+0]),
      .S1 (ConfigBits[372+1]),
      .S1N(ConfigBits_N[372+1]),
      .S2 (ConfigBits[372+2]),
      .S2N(ConfigBits_N[372+2]),
      .S3 (ConfigBits[372+3]),
      .S3N(ConfigBits_N[372+3]),
      .X  (JW2BEG6)
  );

  // switch matrix multiplexer  JW2BEG7         MUX-16
  assign JW2BEG7_input = {
    BD2,
    BD1,
    BD0,
    AD3,
    AD2,
    AD1,
    AD0,
    WW4END0,
    W1END0,
    S2END0,
    S1END2,
    S1END0,
    E2END0,
    E1END0,
    N2END0,
    N1END0
  };
  cus_mux161_buf inst_cus_mux161_buf_JW2BEG7 (
      .A0 (JW2BEG7_input[0]),
      .A1 (JW2BEG7_input[1]),
      .A2 (JW2BEG7_input[2]),
      .A3 (JW2BEG7_input[3]),
      .A4 (JW2BEG7_input[4]),
      .A5 (JW2BEG7_input[5]),
      .A6 (JW2BEG7_input[6]),
      .A7 (JW2BEG7_input[7]),
      .A8 (JW2BEG7_input[8]),
      .A9 (JW2BEG7_input[9]),
      .A10(JW2BEG7_input[10]),
      .A11(JW2BEG7_input[11]),
      .A12(JW2BEG7_input[12]),
      .A13(JW2BEG7_input[13]),
      .A14(JW2BEG7_input[14]),
      .A15(JW2BEG7_input[15]),
      .S0 (ConfigBits[376+0]),
      .S0N(ConfigBits_N[376+0]),
      .S1 (ConfigBits[376+1]),
      .S1N(ConfigBits_N[376+1]),
      .S2 (ConfigBits[376+2]),
      .S2N(ConfigBits_N[376+2]),
      .S3 (ConfigBits[376+3]),
      .S3N(ConfigBits_N[376+3]),
      .X  (JW2BEG7)
  );

  // switch matrix multiplexer  J_l_AB_BEG0         MUX-4
  assign J_l_AB_BEG0_input = {JN2END1, W2END3, S4END3, N4END3};
  cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG0 (
      .A0 (J_l_AB_BEG0_input[0]),
      .A1 (J_l_AB_BEG0_input[1]),
      .A2 (J_l_AB_BEG0_input[2]),
      .A3 (J_l_AB_BEG0_input[3]),
      .S0 (ConfigBits[380+0]),
      .S0N(ConfigBits_N[380+0]),
      .S1 (ConfigBits[380+1]),
      .S1N(ConfigBits_N[380+1]),
      .X  (J_l_AB_BEG0)
  );

  // switch matrix multiplexer  J_l_AB_BEG1         MUX-4
  assign J_l_AB_BEG1_input = {JE2END1, W2END7, S4END2, E2END2};
  cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG1 (
      .A0 (J_l_AB_BEG1_input[0]),
      .A1 (J_l_AB_BEG1_input[1]),
      .A2 (J_l_AB_BEG1_input[2]),
      .A3 (J_l_AB_BEG1_input[3]),
      .S0 (ConfigBits[382+0]),
      .S0N(ConfigBits_N[382+0]),
      .S1 (ConfigBits[382+1]),
      .S1N(ConfigBits_N[382+1]),
      .X  (J_l_AB_BEG1)
  );

  // switch matrix multiplexer  J_l_AB_BEG2         MUX-4
  assign J_l_AB_BEG2_input = {JS2END1, W6END1, E6END1, N4END1};
  cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG2 (
      .A0 (J_l_AB_BEG2_input[0]),
      .A1 (J_l_AB_BEG2_input[1]),
      .A2 (J_l_AB_BEG2_input[2]),
      .A3 (J_l_AB_BEG2_input[3]),
      .S0 (ConfigBits[384+0]),
      .S0N(ConfigBits_N[384+0]),
      .S1 (ConfigBits[384+1]),
      .S1N(ConfigBits_N[384+1]),
      .X  (J_l_AB_BEG2)
  );

  // switch matrix multiplexer  J_l_AB_BEG3         MUX-4
  assign J_l_AB_BEG3_input = {JW2END1, S4END0, E6END0, N4END0};
  cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG3 (
      .A0 (J_l_AB_BEG3_input[0]),
      .A1 (J_l_AB_BEG3_input[1]),
      .A2 (J_l_AB_BEG3_input[2]),
      .A3 (J_l_AB_BEG3_input[3]),
      .S0 (ConfigBits[386+0]),
      .S0N(ConfigBits_N[386+0]),
      .S1 (ConfigBits[386+1]),
      .S1N(ConfigBits_N[386+1]),
      .X  (J_l_AB_BEG3)
  );

  // switch matrix multiplexer  J_l_CD_BEG0         MUX-4
  assign J_l_CD_BEG0_input = {JN2END2, W2END3, S4END3, E2END3};
  cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG0 (
      .A0 (J_l_CD_BEG0_input[0]),
      .A1 (J_l_CD_BEG0_input[1]),
      .A2 (J_l_CD_BEG0_input[2]),
      .A3 (J_l_CD_BEG0_input[3]),
      .S0 (ConfigBits[388+0]),
      .S0N(ConfigBits_N[388+0]),
      .S1 (ConfigBits[388+1]),
      .S1N(ConfigBits_N[388+1]),
      .X  (J_l_CD_BEG0)
  );

  // switch matrix multiplexer  J_l_CD_BEG1         MUX-4
  assign J_l_CD_BEG1_input = {JE2END2, W2END7, E2END2, N4END2};
  cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG1 (
      .A0 (J_l_CD_BEG1_input[0]),
      .A1 (J_l_CD_BEG1_input[1]),
      .A2 (J_l_CD_BEG1_input[2]),
      .A3 (J_l_CD_BEG1_input[3]),
      .S0 (ConfigBits[390+0]),
      .S0N(ConfigBits_N[390+0]),
      .S1 (ConfigBits[390+1]),
      .S1N(ConfigBits_N[390+1]),
      .X  (J_l_CD_BEG1)
  );

  // switch matrix multiplexer  J_l_CD_BEG2         MUX-4
  assign J_l_CD_BEG2_input = {JS2END2, S4END1, E6END1, N4END1};
  cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG2 (
      .A0 (J_l_CD_BEG2_input[0]),
      .A1 (J_l_CD_BEG2_input[1]),
      .A2 (J_l_CD_BEG2_input[2]),
      .A3 (J_l_CD_BEG2_input[3]),
      .S0 (ConfigBits[392+0]),
      .S0N(ConfigBits_N[392+0]),
      .S1 (ConfigBits[392+1]),
      .S1N(ConfigBits_N[392+1]),
      .X  (J_l_CD_BEG2)
  );

  // switch matrix multiplexer  J_l_CD_BEG3         MUX-4
  assign J_l_CD_BEG3_input = {JW2END2, W6END0, S4END0, N4END0};
  cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG3 (
      .A0 (J_l_CD_BEG3_input[0]),
      .A1 (J_l_CD_BEG3_input[1]),
      .A2 (J_l_CD_BEG3_input[2]),
      .A3 (J_l_CD_BEG3_input[3]),
      .S0 (ConfigBits[394+0]),
      .S0N(ConfigBits_N[394+0]),
      .S1 (ConfigBits[394+1]),
      .S1N(ConfigBits_N[394+1]),
      .X  (J_l_CD_BEG3)
  );

  // switch matrix multiplexer  J_l_EF_BEG0         MUX-4
  assign J_l_EF_BEG0_input = {JN2END3, W2END3, E2END3, N4END3};
  cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG0 (
      .A0 (J_l_EF_BEG0_input[0]),
      .A1 (J_l_EF_BEG0_input[1]),
      .A2 (J_l_EF_BEG0_input[2]),
      .A3 (J_l_EF_BEG0_input[3]),
      .S0 (ConfigBits[396+0]),
      .S0N(ConfigBits_N[396+0]),
      .S1 (ConfigBits[396+1]),
      .S1N(ConfigBits_N[396+1]),
      .X  (J_l_EF_BEG0)
  );

  // switch matrix multiplexer  J_l_EF_BEG1         MUX-4
  assign J_l_EF_BEG1_input = {JE2END3, S4END2, E2END2, N4END2};
  cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG1 (
      .A0 (J_l_EF_BEG1_input[0]),
      .A1 (J_l_EF_BEG1_input[1]),
      .A2 (J_l_EF_BEG1_input[2]),
      .A3 (J_l_EF_BEG1_input[3]),
      .S0 (ConfigBits[398+0]),
      .S0N(ConfigBits_N[398+0]),
      .S1 (ConfigBits[398+1]),
      .S1N(ConfigBits_N[398+1]),
      .X  (J_l_EF_BEG1)
  );

  // switch matrix multiplexer  J_l_EF_BEG2         MUX-4
  assign J_l_EF_BEG2_input = {JS2END3, W2END4, S4END1, N4END1};
  cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG2 (
      .A0 (J_l_EF_BEG2_input[0]),
      .A1 (J_l_EF_BEG2_input[1]),
      .A2 (J_l_EF_BEG2_input[2]),
      .A3 (J_l_EF_BEG2_input[3]),
      .S0 (ConfigBits[400+0]),
      .S0N(ConfigBits_N[400+0]),
      .S1 (ConfigBits[400+1]),
      .S1N(ConfigBits_N[400+1]),
      .X  (J_l_EF_BEG2)
  );

  // switch matrix multiplexer  J_l_EF_BEG3         MUX-4
  assign J_l_EF_BEG3_input = {JW2END3, W2END0, S4END0, E6END0};
  cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG3 (
      .A0 (J_l_EF_BEG3_input[0]),
      .A1 (J_l_EF_BEG3_input[1]),
      .A2 (J_l_EF_BEG3_input[2]),
      .A3 (J_l_EF_BEG3_input[3]),
      .S0 (ConfigBits[402+0]),
      .S0N(ConfigBits_N[402+0]),
      .S1 (ConfigBits[402+1]),
      .S1N(ConfigBits_N[402+1]),
      .X  (J_l_EF_BEG3)
  );

  // switch matrix multiplexer  J_l_GH_BEG0         MUX-4
  assign J_l_GH_BEG0_input = {JN2END4, S4END3, E2END3, N4END3};
  cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG0 (
      .A0 (J_l_GH_BEG0_input[0]),
      .A1 (J_l_GH_BEG0_input[1]),
      .A2 (J_l_GH_BEG0_input[2]),
      .A3 (J_l_GH_BEG0_input[3]),
      .S0 (ConfigBits[404+0]),
      .S0N(ConfigBits_N[404+0]),
      .S1 (ConfigBits[404+1]),
      .S1N(ConfigBits_N[404+1]),
      .X  (J_l_GH_BEG0)
  );

  // switch matrix multiplexer  J_l_GH_BEG1         MUX-4
  assign J_l_GH_BEG1_input = {JE2END4, W2END2, S4END2, N4END2};
  cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG1 (
      .A0 (J_l_GH_BEG1_input[0]),
      .A1 (J_l_GH_BEG1_input[1]),
      .A2 (J_l_GH_BEG1_input[2]),
      .A3 (J_l_GH_BEG1_input[3]),
      .S0 (ConfigBits[406+0]),
      .S0N(ConfigBits_N[406+0]),
      .S1 (ConfigBits[406+1]),
      .S1N(ConfigBits_N[406+1]),
      .X  (J_l_GH_BEG1)
  );

  // switch matrix multiplexer  J_l_GH_BEG2         MUX-4
  assign J_l_GH_BEG2_input = {JS2END4, W2END4, S4END1, E6END1};
  cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG2 (
      .A0 (J_l_GH_BEG2_input[0]),
      .A1 (J_l_GH_BEG2_input[1]),
      .A2 (J_l_GH_BEG2_input[2]),
      .A3 (J_l_GH_BEG2_input[3]),
      .S0 (ConfigBits[408+0]),
      .S0N(ConfigBits_N[408+0]),
      .S1 (ConfigBits[408+1]),
      .S1N(ConfigBits_N[408+1]),
      .X  (J_l_GH_BEG2)
  );

  // switch matrix multiplexer  J_l_GH_BEG3         MUX-4
  assign J_l_GH_BEG3_input = {JW2END4, W2END0, E6END0, N4END0};
  cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG3 (
      .A0 (J_l_GH_BEG3_input[0]),
      .A1 (J_l_GH_BEG3_input[1]),
      .A2 (J_l_GH_BEG3_input[2]),
      .A3 (J_l_GH_BEG3_input[3]),
      .S0 (ConfigBits[410+0]),
      .S0N(ConfigBits_N[410+0]),
      .S1 (ConfigBits[410+1]),
      .S1N(ConfigBits_N[410+1]),
      .X  (J_l_GH_BEG3)
  );

  assign DEBUG_select_N1BEG0 = ConfigBits[1:0];
  assign DEBUG_select_N1BEG1 = ConfigBits[3:2];
  assign DEBUG_select_N1BEG2 = ConfigBits[5:4];
  assign DEBUG_select_N1BEG3 = ConfigBits[7:6];
  assign DEBUG_select_N4BEG0 = ConfigBits[9:8];
  assign DEBUG_select_N4BEG1 = ConfigBits[11:10];
  assign DEBUG_select_N4BEG2 = ConfigBits[13:12];
  assign DEBUG_select_N4BEG3 = ConfigBits[15:14];
  assign DEBUG_select_NN4BEG0 = ConfigBits[18:16];
  assign DEBUG_select_NN4BEG1 = ConfigBits[21:19];
  assign DEBUG_select_NN4BEG2 = ConfigBits[24:22];
  assign DEBUG_select_NN4BEG3 = ConfigBits[27:25];
  assign DEBUG_select_E1BEG0 = ConfigBits[29:28];
  assign DEBUG_select_E1BEG1 = ConfigBits[31:30];
  assign DEBUG_select_E1BEG2 = ConfigBits[33:32];
  assign DEBUG_select_E1BEG3 = ConfigBits[35:34];
  assign DEBUG_select_EE4BEG0 = ConfigBits[38:36];
  assign DEBUG_select_EE4BEG1 = ConfigBits[41:39];
  assign DEBUG_select_EE4BEG2 = ConfigBits[44:42];
  assign DEBUG_select_EE4BEG3 = ConfigBits[47:45];
  assign DEBUG_select_E6BEG0 = ConfigBits[51:48];
  assign DEBUG_select_E6BEG1 = ConfigBits[55:52];
  assign DEBUG_select_S1BEG0 = ConfigBits[57:56];
  assign DEBUG_select_S1BEG1 = ConfigBits[59:58];
  assign DEBUG_select_S1BEG2 = ConfigBits[61:60];
  assign DEBUG_select_S1BEG3 = ConfigBits[63:62];
  assign DEBUG_select_S4BEG0 = ConfigBits[65:64];
  assign DEBUG_select_S4BEG1 = ConfigBits[67:66];
  assign DEBUG_select_S4BEG2 = ConfigBits[69:68];
  assign DEBUG_select_S4BEG3 = ConfigBits[71:70];
  assign DEBUG_select_SS4BEG0 = ConfigBits[74:72];
  assign DEBUG_select_SS4BEG1 = ConfigBits[77:75];
  assign DEBUG_select_SS4BEG2 = ConfigBits[80:78];
  assign DEBUG_select_SS4BEG3 = ConfigBits[83:81];
  assign DEBUG_select_W1BEG0 = ConfigBits[85:84];
  assign DEBUG_select_W1BEG1 = ConfigBits[87:86];
  assign DEBUG_select_W1BEG2 = ConfigBits[89:88];
  assign DEBUG_select_W1BEG3 = ConfigBits[91:90];
  assign DEBUG_select_WW4BEG0 = ConfigBits[94:92];
  assign DEBUG_select_WW4BEG1 = ConfigBits[97:95];
  assign DEBUG_select_WW4BEG2 = ConfigBits[100:98];
  assign DEBUG_select_WW4BEG3 = ConfigBits[103:101];
  assign DEBUG_select_W6BEG0 = ConfigBits[107:104];
  assign DEBUG_select_W6BEG1 = ConfigBits[111:108];
  assign DEBUG_select_D0 = ConfigBits[113:112];
  assign DEBUG_select_D1 = ConfigBits[115:114];
  assign DEBUG_select_D2 = ConfigBits[117:116];
  assign DEBUG_select_D3 = ConfigBits[119:118];
  assign DEBUG_select_W_ADR0 = ConfigBits[121:120];
  assign DEBUG_select_W_ADR1 = ConfigBits[123:122];
  assign DEBUG_select_W_ADR2 = ConfigBits[125:124];
  assign DEBUG_select_W_ADR3 = ConfigBits[127:126];
  assign DEBUG_select_W_ADR4 = ConfigBits[130:128];
  assign DEBUG_select_W_en = ConfigBits[133:131];
  assign DEBUG_select_A_ADR0 = ConfigBits[135:134];
  assign DEBUG_select_A_ADR1 = ConfigBits[137:136];
  assign DEBUG_select_A_ADR2 = ConfigBits[139:138];
  assign DEBUG_select_A_ADR3 = ConfigBits[141:140];
  assign DEBUG_select_A_ADR4 = ConfigBits[144:142];
  assign DEBUG_select_B_ADR0 = ConfigBits[146:145];
  assign DEBUG_select_B_ADR1 = ConfigBits[148:147];
  assign DEBUG_select_B_ADR2 = ConfigBits[150:149];
  assign DEBUG_select_B_ADR3 = ConfigBits[152:151];
  assign DEBUG_select_B_ADR4 = ConfigBits[155:153];
  assign DEBUG_select_J2MID_ABa_BEG0 = ConfigBits[157:156];
  assign DEBUG_select_J2MID_ABa_BEG1 = ConfigBits[159:158];
  assign DEBUG_select_J2MID_ABa_BEG2 = ConfigBits[161:160];
  assign DEBUG_select_J2MID_ABa_BEG3 = ConfigBits[163:162];
  assign DEBUG_select_J2MID_CDa_BEG0 = ConfigBits[165:164];
  assign DEBUG_select_J2MID_CDa_BEG1 = ConfigBits[167:166];
  assign DEBUG_select_J2MID_CDa_BEG2 = ConfigBits[169:168];
  assign DEBUG_select_J2MID_CDa_BEG3 = ConfigBits[171:170];
  assign DEBUG_select_J2MID_EFa_BEG0 = ConfigBits[173:172];
  assign DEBUG_select_J2MID_EFa_BEG1 = ConfigBits[175:174];
  assign DEBUG_select_J2MID_EFa_BEG2 = ConfigBits[177:176];
  assign DEBUG_select_J2MID_EFa_BEG3 = ConfigBits[179:178];
  assign DEBUG_select_J2MID_GHa_BEG0 = ConfigBits[181:180];
  assign DEBUG_select_J2MID_GHa_BEG1 = ConfigBits[183:182];
  assign DEBUG_select_J2MID_GHa_BEG2 = ConfigBits[185:184];
  assign DEBUG_select_J2MID_GHa_BEG3 = ConfigBits[187:186];
  assign DEBUG_select_J2MID_ABb_BEG0 = ConfigBits[189:188];
  assign DEBUG_select_J2MID_ABb_BEG1 = ConfigBits[191:190];
  assign DEBUG_select_J2MID_ABb_BEG2 = ConfigBits[193:192];
  assign DEBUG_select_J2MID_ABb_BEG3 = ConfigBits[195:194];
  assign DEBUG_select_J2MID_CDb_BEG0 = ConfigBits[197:196];
  assign DEBUG_select_J2MID_CDb_BEG1 = ConfigBits[199:198];
  assign DEBUG_select_J2MID_CDb_BEG2 = ConfigBits[201:200];
  assign DEBUG_select_J2MID_CDb_BEG3 = ConfigBits[203:202];
  assign DEBUG_select_J2MID_EFb_BEG0 = ConfigBits[205:204];
  assign DEBUG_select_J2MID_EFb_BEG1 = ConfigBits[207:206];
  assign DEBUG_select_J2MID_EFb_BEG2 = ConfigBits[209:208];
  assign DEBUG_select_J2MID_EFb_BEG3 = ConfigBits[211:210];
  assign DEBUG_select_J2MID_GHb_BEG0 = ConfigBits[213:212];
  assign DEBUG_select_J2MID_GHb_BEG1 = ConfigBits[215:214];
  assign DEBUG_select_J2MID_GHb_BEG2 = ConfigBits[217:216];
  assign DEBUG_select_J2MID_GHb_BEG3 = ConfigBits[219:218];
  assign DEBUG_select_J2END_AB_BEG0 = ConfigBits[221:220];
  assign DEBUG_select_J2END_AB_BEG1 = ConfigBits[223:222];
  assign DEBUG_select_J2END_AB_BEG2 = ConfigBits[225:224];
  assign DEBUG_select_J2END_AB_BEG3 = ConfigBits[227:226];
  assign DEBUG_select_J2END_CD_BEG0 = ConfigBits[229:228];
  assign DEBUG_select_J2END_CD_BEG1 = ConfigBits[231:230];
  assign DEBUG_select_J2END_CD_BEG2 = ConfigBits[233:232];
  assign DEBUG_select_J2END_CD_BEG3 = ConfigBits[235:234];
  assign DEBUG_select_J2END_EF_BEG0 = ConfigBits[237:236];
  assign DEBUG_select_J2END_EF_BEG1 = ConfigBits[239:238];
  assign DEBUG_select_J2END_EF_BEG2 = ConfigBits[241:240];
  assign DEBUG_select_J2END_EF_BEG3 = ConfigBits[243:242];
  assign DEBUG_select_J2END_GH_BEG0 = ConfigBits[245:244];
  assign DEBUG_select_J2END_GH_BEG1 = ConfigBits[247:246];
  assign DEBUG_select_J2END_GH_BEG2 = ConfigBits[249:248];
  assign DEBUG_select_J2END_GH_BEG3 = ConfigBits[251:250];
  assign DEBUG_select_JN2BEG0 = ConfigBits[255:252];
  assign DEBUG_select_JN2BEG1 = ConfigBits[259:256];
  assign DEBUG_select_JN2BEG2 = ConfigBits[263:260];
  assign DEBUG_select_JN2BEG3 = ConfigBits[267:264];
  assign DEBUG_select_JN2BEG4 = ConfigBits[271:268];
  assign DEBUG_select_JN2BEG5 = ConfigBits[275:272];
  assign DEBUG_select_JN2BEG6 = ConfigBits[279:276];
  assign DEBUG_select_JN2BEG7 = ConfigBits[283:280];
  assign DEBUG_select_JE2BEG0 = ConfigBits[287:284];
  assign DEBUG_select_JE2BEG1 = ConfigBits[291:288];
  assign DEBUG_select_JE2BEG2 = ConfigBits[295:292];
  assign DEBUG_select_JE2BEG3 = ConfigBits[299:296];
  assign DEBUG_select_JE2BEG4 = ConfigBits[303:300];
  assign DEBUG_select_JE2BEG5 = ConfigBits[307:304];
  assign DEBUG_select_JE2BEG6 = ConfigBits[311:308];
  assign DEBUG_select_JE2BEG7 = ConfigBits[315:312];
  assign DEBUG_select_JS2BEG0 = ConfigBits[319:316];
  assign DEBUG_select_JS2BEG1 = ConfigBits[323:320];
  assign DEBUG_select_JS2BEG2 = ConfigBits[327:324];
  assign DEBUG_select_JS2BEG3 = ConfigBits[331:328];
  assign DEBUG_select_JS2BEG4 = ConfigBits[335:332];
  assign DEBUG_select_JS2BEG5 = ConfigBits[339:336];
  assign DEBUG_select_JS2BEG6 = ConfigBits[343:340];
  assign DEBUG_select_JS2BEG7 = ConfigBits[347:344];
  assign DEBUG_select_JW2BEG0 = ConfigBits[351:348];
  assign DEBUG_select_JW2BEG1 = ConfigBits[355:352];
  assign DEBUG_select_JW2BEG2 = ConfigBits[359:356];
  assign DEBUG_select_JW2BEG3 = ConfigBits[363:360];
  assign DEBUG_select_JW2BEG4 = ConfigBits[367:364];
  assign DEBUG_select_JW2BEG5 = ConfigBits[371:368];
  assign DEBUG_select_JW2BEG6 = ConfigBits[375:372];
  assign DEBUG_select_JW2BEG7 = ConfigBits[379:376];
  assign DEBUG_select_J_l_AB_BEG0 = ConfigBits[381:380];
  assign DEBUG_select_J_l_AB_BEG1 = ConfigBits[383:382];
  assign DEBUG_select_J_l_AB_BEG2 = ConfigBits[385:384];
  assign DEBUG_select_J_l_AB_BEG3 = ConfigBits[387:386];
  assign DEBUG_select_J_l_CD_BEG0 = ConfigBits[389:388];
  assign DEBUG_select_J_l_CD_BEG1 = ConfigBits[391:390];
  assign DEBUG_select_J_l_CD_BEG2 = ConfigBits[393:392];
  assign DEBUG_select_J_l_CD_BEG3 = ConfigBits[395:394];
  assign DEBUG_select_J_l_EF_BEG0 = ConfigBits[397:396];
  assign DEBUG_select_J_l_EF_BEG1 = ConfigBits[399:398];
  assign DEBUG_select_J_l_EF_BEG2 = ConfigBits[401:400];
  assign DEBUG_select_J_l_EF_BEG3 = ConfigBits[403:402];
  assign DEBUG_select_J_l_GH_BEG0 = ConfigBits[405:404];
  assign DEBUG_select_J_l_GH_BEG1 = ConfigBits[407:406];
  assign DEBUG_select_J_l_GH_BEG2 = ConfigBits[409:408];
  assign DEBUG_select_J_l_GH_BEG3 = ConfigBits[411:410];

endmodule
